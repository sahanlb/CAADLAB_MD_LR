localparam [GSIZE1DX-1:0][GSIZE1DY-1:0][GSIZE1DZ-1:0][1:0][31:0] GMEM_IFFTY_CHK = {
  {32'h43adb08f, 32'hc36eab13} /* (31, 31, 31) {real, imag} */,
  {32'hc38c81aa, 32'h4341a2f8} /* (31, 31, 30) {real, imag} */,
  {32'h3ff2d970, 32'hc1ae82e6} /* (31, 31, 29) {real, imag} */,
  {32'h428aba9c, 32'h425dba23} /* (31, 31, 28) {real, imag} */,
  {32'hc26ff125, 32'h419abe34} /* (31, 31, 27) {real, imag} */,
  {32'h3ff629c0, 32'hc1497c9a} /* (31, 31, 26) {real, imag} */,
  {32'hc19bfc9a, 32'hc1f6848a} /* (31, 31, 25) {real, imag} */,
  {32'h420a7628, 32'h423ee6ee} /* (31, 31, 24) {real, imag} */,
  {32'hc214d280, 32'h419852e5} /* (31, 31, 23) {real, imag} */,
  {32'hc196cedb, 32'hc20fbaf3} /* (31, 31, 22) {real, imag} */,
  {32'hc20cd3d0, 32'h4176c7cd} /* (31, 31, 21) {real, imag} */,
  {32'h421f948c, 32'hc212eb88} /* (31, 31, 20) {real, imag} */,
  {32'h419101b8, 32'h415684b1} /* (31, 31, 19) {real, imag} */,
  {32'h41df04c4, 32'hbfb3c2c8} /* (31, 31, 18) {real, imag} */,
  {32'h4183bb16, 32'hc17b7f98} /* (31, 31, 17) {real, imag} */,
  {32'hc0233e80, 32'h00000000} /* (31, 31, 16) {real, imag} */,
  {32'h4183bb16, 32'h417b7f98} /* (31, 31, 15) {real, imag} */,
  {32'h41df04c4, 32'h3fb3c2c8} /* (31, 31, 14) {real, imag} */,
  {32'h419101b8, 32'hc15684b1} /* (31, 31, 13) {real, imag} */,
  {32'h421f948c, 32'h4212eb88} /* (31, 31, 12) {real, imag} */,
  {32'hc20cd3d0, 32'hc176c7cd} /* (31, 31, 11) {real, imag} */,
  {32'hc196cedb, 32'h420fbaf3} /* (31, 31, 10) {real, imag} */,
  {32'hc214d280, 32'hc19852e5} /* (31, 31, 9) {real, imag} */,
  {32'h420a7628, 32'hc23ee6ee} /* (31, 31, 8) {real, imag} */,
  {32'hc19bfc9a, 32'h41f6848a} /* (31, 31, 7) {real, imag} */,
  {32'h3ff629c0, 32'h41497c9a} /* (31, 31, 6) {real, imag} */,
  {32'hc26ff125, 32'hc19abe34} /* (31, 31, 5) {real, imag} */,
  {32'h428aba9c, 32'hc25dba23} /* (31, 31, 4) {real, imag} */,
  {32'h3ff2d970, 32'h41ae82e6} /* (31, 31, 3) {real, imag} */,
  {32'hc38c81aa, 32'hc341a2f8} /* (31, 31, 2) {real, imag} */,
  {32'h43adb08f, 32'h436eab13} /* (31, 31, 1) {real, imag} */,
  {32'h4361b5c3, 32'h00000000} /* (31, 31, 0) {real, imag} */,
  {32'h4406c004, 32'hc38db278} /* (31, 30, 31) {real, imag} */,
  {32'hc3e68306, 32'h438c601a} /* (31, 30, 30) {real, imag} */,
  {32'h41a503bc, 32'hbe6cf200} /* (31, 30, 29) {real, imag} */,
  {32'h4260a8d2, 32'h3f848b00} /* (31, 30, 28) {real, imag} */,
  {32'hc2331a3b, 32'h41b4e6eb} /* (31, 30, 27) {real, imag} */,
  {32'h42298a0a, 32'hbfdc6040} /* (31, 30, 26) {real, imag} */,
  {32'hc20da2f1, 32'hc2a17a32} /* (31, 30, 25) {real, imag} */,
  {32'h429fd303, 32'h41fa05ce} /* (31, 30, 24) {real, imag} */,
  {32'hc028fc40, 32'hc280b69a} /* (31, 30, 23) {real, imag} */,
  {32'hc27098d0, 32'hbfb30bc0} /* (31, 30, 22) {real, imag} */,
  {32'hc21ca92a, 32'hc05135a4} /* (31, 30, 21) {real, imag} */,
  {32'h403b81e0, 32'hc1a89e92} /* (31, 30, 20) {real, imag} */,
  {32'h4118aed2, 32'h40357140} /* (31, 30, 19) {real, imag} */,
  {32'h428c26ba, 32'hc13db234} /* (31, 30, 18) {real, imag} */,
  {32'hc190fae4, 32'hc0e51205} /* (31, 30, 17) {real, imag} */,
  {32'hc21e14e9, 32'h00000000} /* (31, 30, 16) {real, imag} */,
  {32'hc190fae4, 32'h40e51205} /* (31, 30, 15) {real, imag} */,
  {32'h428c26ba, 32'h413db234} /* (31, 30, 14) {real, imag} */,
  {32'h4118aed2, 32'hc0357140} /* (31, 30, 13) {real, imag} */,
  {32'h403b81e0, 32'h41a89e92} /* (31, 30, 12) {real, imag} */,
  {32'hc21ca92a, 32'h405135a4} /* (31, 30, 11) {real, imag} */,
  {32'hc27098d0, 32'h3fb30bc0} /* (31, 30, 10) {real, imag} */,
  {32'hc028fc40, 32'h4280b69a} /* (31, 30, 9) {real, imag} */,
  {32'h429fd303, 32'hc1fa05ce} /* (31, 30, 8) {real, imag} */,
  {32'hc20da2f1, 32'h42a17a32} /* (31, 30, 7) {real, imag} */,
  {32'h42298a0a, 32'h3fdc6040} /* (31, 30, 6) {real, imag} */,
  {32'hc2331a3b, 32'hc1b4e6eb} /* (31, 30, 5) {real, imag} */,
  {32'h4260a8d2, 32'hbf848b00} /* (31, 30, 4) {real, imag} */,
  {32'h41a503bc, 32'h3e6cf200} /* (31, 30, 3) {real, imag} */,
  {32'hc3e68306, 32'hc38c601a} /* (31, 30, 2) {real, imag} */,
  {32'h4406c004, 32'h438db278} /* (31, 30, 1) {real, imag} */,
  {32'h433a5132, 32'h00000000} /* (31, 30, 0) {real, imag} */,
  {32'h441ba38e, 32'hc3207cd1} /* (31, 29, 31) {real, imag} */,
  {32'hc3c2b284, 32'h437a9433} /* (31, 29, 30) {real, imag} */,
  {32'hc15e4818, 32'h42905a4f} /* (31, 29, 29) {real, imag} */,
  {32'h42c1f415, 32'h40aaa560} /* (31, 29, 28) {real, imag} */,
  {32'hc280f407, 32'h41636fac} /* (31, 29, 27) {real, imag} */,
  {32'hc2821fcc, 32'hc1a91dcc} /* (31, 29, 26) {real, imag} */,
  {32'h418d592e, 32'hc20a6626} /* (31, 29, 25) {real, imag} */,
  {32'hc1f2439b, 32'h41bf5be2} /* (31, 29, 24) {real, imag} */,
  {32'hc1475fa7, 32'h42d6ceb8} /* (31, 29, 23) {real, imag} */,
  {32'h4276be28, 32'hc2270a68} /* (31, 29, 22) {real, imag} */,
  {32'hc252fb64, 32'hc1f4fea7} /* (31, 29, 21) {real, imag} */,
  {32'hc19ac18a, 32'h422c1d84} /* (31, 29, 20) {real, imag} */,
  {32'hbfc447c0, 32'hc2ece47f} /* (31, 29, 19) {real, imag} */,
  {32'hc1b0ba27, 32'hc1faf237} /* (31, 29, 18) {real, imag} */,
  {32'hc1ba963a, 32'hc1ad5670} /* (31, 29, 17) {real, imag} */,
  {32'h4293ec56, 32'h00000000} /* (31, 29, 16) {real, imag} */,
  {32'hc1ba963a, 32'h41ad5670} /* (31, 29, 15) {real, imag} */,
  {32'hc1b0ba27, 32'h41faf237} /* (31, 29, 14) {real, imag} */,
  {32'hbfc447c0, 32'h42ece47f} /* (31, 29, 13) {real, imag} */,
  {32'hc19ac18a, 32'hc22c1d84} /* (31, 29, 12) {real, imag} */,
  {32'hc252fb64, 32'h41f4fea7} /* (31, 29, 11) {real, imag} */,
  {32'h4276be28, 32'h42270a68} /* (31, 29, 10) {real, imag} */,
  {32'hc1475fa7, 32'hc2d6ceb8} /* (31, 29, 9) {real, imag} */,
  {32'hc1f2439b, 32'hc1bf5be2} /* (31, 29, 8) {real, imag} */,
  {32'h418d592e, 32'h420a6626} /* (31, 29, 7) {real, imag} */,
  {32'hc2821fcc, 32'h41a91dcc} /* (31, 29, 6) {real, imag} */,
  {32'hc280f407, 32'hc1636fac} /* (31, 29, 5) {real, imag} */,
  {32'h42c1f415, 32'hc0aaa560} /* (31, 29, 4) {real, imag} */,
  {32'hc15e4818, 32'hc2905a4f} /* (31, 29, 3) {real, imag} */,
  {32'hc3c2b284, 32'hc37a9433} /* (31, 29, 2) {real, imag} */,
  {32'h441ba38e, 32'h43207cd1} /* (31, 29, 1) {real, imag} */,
  {32'h43389a35, 32'h00000000} /* (31, 29, 0) {real, imag} */,
  {32'h440b6094, 32'hc2e882c6} /* (31, 28, 31) {real, imag} */,
  {32'hc396625b, 32'h42b48b90} /* (31, 28, 30) {real, imag} */,
  {32'hc2237ab7, 32'hc0e41b3e} /* (31, 28, 29) {real, imag} */,
  {32'h431d85c8, 32'h427a02c5} /* (31, 28, 28) {real, imag} */,
  {32'hc297176f, 32'hc1edfe16} /* (31, 28, 27) {real, imag} */,
  {32'hc178ccc0, 32'h4296b304} /* (31, 28, 26) {real, imag} */,
  {32'h40de2dc4, 32'hc2878784} /* (31, 28, 25) {real, imag} */,
  {32'hc2a60d7c, 32'h42c8e82e} /* (31, 28, 24) {real, imag} */,
  {32'h4221c1c9, 32'h41b6de37} /* (31, 28, 23) {real, imag} */,
  {32'hc13c8226, 32'hc145ff2b} /* (31, 28, 22) {real, imag} */,
  {32'hc178758f, 32'hc194a35e} /* (31, 28, 21) {real, imag} */,
  {32'h40f6a138, 32'hc1b7484a} /* (31, 28, 20) {real, imag} */,
  {32'hc14c789f, 32'h420a334f} /* (31, 28, 19) {real, imag} */,
  {32'hc22b79ca, 32'h425a84ef} /* (31, 28, 18) {real, imag} */,
  {32'h4230f1f1, 32'hc0fa8b83} /* (31, 28, 17) {real, imag} */,
  {32'hc1075eae, 32'h00000000} /* (31, 28, 16) {real, imag} */,
  {32'h4230f1f1, 32'h40fa8b83} /* (31, 28, 15) {real, imag} */,
  {32'hc22b79ca, 32'hc25a84ef} /* (31, 28, 14) {real, imag} */,
  {32'hc14c789f, 32'hc20a334f} /* (31, 28, 13) {real, imag} */,
  {32'h40f6a138, 32'h41b7484a} /* (31, 28, 12) {real, imag} */,
  {32'hc178758f, 32'h4194a35e} /* (31, 28, 11) {real, imag} */,
  {32'hc13c8226, 32'h4145ff2b} /* (31, 28, 10) {real, imag} */,
  {32'h4221c1c9, 32'hc1b6de37} /* (31, 28, 9) {real, imag} */,
  {32'hc2a60d7c, 32'hc2c8e82e} /* (31, 28, 8) {real, imag} */,
  {32'h40de2dc4, 32'h42878784} /* (31, 28, 7) {real, imag} */,
  {32'hc178ccc0, 32'hc296b304} /* (31, 28, 6) {real, imag} */,
  {32'hc297176f, 32'h41edfe16} /* (31, 28, 5) {real, imag} */,
  {32'h431d85c8, 32'hc27a02c5} /* (31, 28, 4) {real, imag} */,
  {32'hc2237ab7, 32'h40e41b3e} /* (31, 28, 3) {real, imag} */,
  {32'hc396625b, 32'hc2b48b90} /* (31, 28, 2) {real, imag} */,
  {32'h440b6094, 32'h42e882c6} /* (31, 28, 1) {real, imag} */,
  {32'h438ddf70, 32'h00000000} /* (31, 28, 0) {real, imag} */,
  {32'h43e36cba, 32'hc30579e5} /* (31, 27, 31) {real, imag} */,
  {32'hc3cc8cdc, 32'h42ffcad0} /* (31, 27, 30) {real, imag} */,
  {32'hc189f400, 32'hc21feb64} /* (31, 27, 29) {real, imag} */,
  {32'hc146aa00, 32'h429e4b84} /* (31, 27, 28) {real, imag} */,
  {32'h4217741e, 32'h40f8dc70} /* (31, 27, 27) {real, imag} */,
  {32'h42094c93, 32'hc1a4344d} /* (31, 27, 26) {real, imag} */,
  {32'hc221dfa4, 32'hc2a19258} /* (31, 27, 25) {real, imag} */,
  {32'hc292d7c7, 32'hc18d0fcd} /* (31, 27, 24) {real, imag} */,
  {32'hbf33c9e0, 32'h421f17a8} /* (31, 27, 23) {real, imag} */,
  {32'h420bf176, 32'hc2227b7e} /* (31, 27, 22) {real, imag} */,
  {32'hc27c6ee2, 32'hbe3a2a00} /* (31, 27, 21) {real, imag} */,
  {32'h41dc435a, 32'h4133fa6e} /* (31, 27, 20) {real, imag} */,
  {32'hc100fde0, 32'h426e8688} /* (31, 27, 19) {real, imag} */,
  {32'hc109948c, 32'h42bfc806} /* (31, 27, 18) {real, imag} */,
  {32'h4197a49e, 32'hc26ceac4} /* (31, 27, 17) {real, imag} */,
  {32'h4223ceaa, 32'h00000000} /* (31, 27, 16) {real, imag} */,
  {32'h4197a49e, 32'h426ceac4} /* (31, 27, 15) {real, imag} */,
  {32'hc109948c, 32'hc2bfc806} /* (31, 27, 14) {real, imag} */,
  {32'hc100fde0, 32'hc26e8688} /* (31, 27, 13) {real, imag} */,
  {32'h41dc435a, 32'hc133fa6e} /* (31, 27, 12) {real, imag} */,
  {32'hc27c6ee2, 32'h3e3a2a00} /* (31, 27, 11) {real, imag} */,
  {32'h420bf176, 32'h42227b7e} /* (31, 27, 10) {real, imag} */,
  {32'hbf33c9e0, 32'hc21f17a8} /* (31, 27, 9) {real, imag} */,
  {32'hc292d7c7, 32'h418d0fcd} /* (31, 27, 8) {real, imag} */,
  {32'hc221dfa4, 32'h42a19258} /* (31, 27, 7) {real, imag} */,
  {32'h42094c93, 32'h41a4344d} /* (31, 27, 6) {real, imag} */,
  {32'h4217741e, 32'hc0f8dc70} /* (31, 27, 5) {real, imag} */,
  {32'hc146aa00, 32'hc29e4b84} /* (31, 27, 4) {real, imag} */,
  {32'hc189f400, 32'h421feb64} /* (31, 27, 3) {real, imag} */,
  {32'hc3cc8cdc, 32'hc2ffcad0} /* (31, 27, 2) {real, imag} */,
  {32'h43e36cba, 32'h430579e5} /* (31, 27, 1) {real, imag} */,
  {32'h43cc18c6, 32'h00000000} /* (31, 27, 0) {real, imag} */,
  {32'h4400b433, 32'hc3151bde} /* (31, 26, 31) {real, imag} */,
  {32'hc403c0fb, 32'h4365101a} /* (31, 26, 30) {real, imag} */,
  {32'h419ca018, 32'hc1549fd9} /* (31, 26, 29) {real, imag} */,
  {32'h420b4f3c, 32'h41cebd44} /* (31, 26, 28) {real, imag} */,
  {32'h4218adee, 32'h41ed3c44} /* (31, 26, 27) {real, imag} */,
  {32'hc1086763, 32'h42153755} /* (31, 26, 26) {real, imag} */,
  {32'hc2461488, 32'hc2aa928a} /* (31, 26, 25) {real, imag} */,
  {32'hc0a32dba, 32'h4253c0e3} /* (31, 26, 24) {real, imag} */,
  {32'hc2b30c44, 32'hc270a386} /* (31, 26, 23) {real, imag} */,
  {32'hc195e595, 32'h4214a8a3} /* (31, 26, 22) {real, imag} */,
  {32'h4213b8fa, 32'h3e6c6200} /* (31, 26, 21) {real, imag} */,
  {32'h41f13308, 32'h421b008c} /* (31, 26, 20) {real, imag} */,
  {32'hc1c2ca25, 32'hc2bfa7e6} /* (31, 26, 19) {real, imag} */,
  {32'hc1be1388, 32'h41f99d08} /* (31, 26, 18) {real, imag} */,
  {32'h4152b2b4, 32'hc1c6f1aa} /* (31, 26, 17) {real, imag} */,
  {32'hc178511b, 32'h00000000} /* (31, 26, 16) {real, imag} */,
  {32'h4152b2b4, 32'h41c6f1aa} /* (31, 26, 15) {real, imag} */,
  {32'hc1be1388, 32'hc1f99d08} /* (31, 26, 14) {real, imag} */,
  {32'hc1c2ca25, 32'h42bfa7e6} /* (31, 26, 13) {real, imag} */,
  {32'h41f13308, 32'hc21b008c} /* (31, 26, 12) {real, imag} */,
  {32'h4213b8fa, 32'hbe6c6200} /* (31, 26, 11) {real, imag} */,
  {32'hc195e595, 32'hc214a8a3} /* (31, 26, 10) {real, imag} */,
  {32'hc2b30c44, 32'h4270a386} /* (31, 26, 9) {real, imag} */,
  {32'hc0a32dba, 32'hc253c0e3} /* (31, 26, 8) {real, imag} */,
  {32'hc2461488, 32'h42aa928a} /* (31, 26, 7) {real, imag} */,
  {32'hc1086763, 32'hc2153755} /* (31, 26, 6) {real, imag} */,
  {32'h4218adee, 32'hc1ed3c44} /* (31, 26, 5) {real, imag} */,
  {32'h420b4f3c, 32'hc1cebd44} /* (31, 26, 4) {real, imag} */,
  {32'h419ca018, 32'h41549fd9} /* (31, 26, 3) {real, imag} */,
  {32'hc403c0fb, 32'hc365101a} /* (31, 26, 2) {real, imag} */,
  {32'h4400b433, 32'h43151bde} /* (31, 26, 1) {real, imag} */,
  {32'h43c8d262, 32'h00000000} /* (31, 26, 0) {real, imag} */,
  {32'h4412f89d, 32'hc13b7963} /* (31, 25, 31) {real, imag} */,
  {32'hc4096ca3, 32'h438b3aea} /* (31, 25, 30) {real, imag} */,
  {32'hc24691f8, 32'h402508e0} /* (31, 25, 29) {real, imag} */,
  {32'h425bea2d, 32'hc23e147a} /* (31, 25, 28) {real, imag} */,
  {32'hc0de0b48, 32'h41e48782} /* (31, 25, 27) {real, imag} */,
  {32'h3fb05340, 32'hc227d4b6} /* (31, 25, 26) {real, imag} */,
  {32'h424db3ea, 32'hc20331d6} /* (31, 25, 25) {real, imag} */,
  {32'hc29a9203, 32'h41b4e7b8} /* (31, 25, 24) {real, imag} */,
  {32'hbe045c00, 32'h4223cc4e} /* (31, 25, 23) {real, imag} */,
  {32'h40b70928, 32'hc17add52} /* (31, 25, 22) {real, imag} */,
  {32'hc2a98860, 32'hc184e68f} /* (31, 25, 21) {real, imag} */,
  {32'h42d318c0, 32'hc1afe4a8} /* (31, 25, 20) {real, imag} */,
  {32'h4286d4b8, 32'hc14049ba} /* (31, 25, 19) {real, imag} */,
  {32'h41a6ea8d, 32'h41a51a27} /* (31, 25, 18) {real, imag} */,
  {32'hc2061826, 32'h429a9658} /* (31, 25, 17) {real, imag} */,
  {32'hc0c1411c, 32'h00000000} /* (31, 25, 16) {real, imag} */,
  {32'hc2061826, 32'hc29a9658} /* (31, 25, 15) {real, imag} */,
  {32'h41a6ea8d, 32'hc1a51a27} /* (31, 25, 14) {real, imag} */,
  {32'h4286d4b8, 32'h414049ba} /* (31, 25, 13) {real, imag} */,
  {32'h42d318c0, 32'h41afe4a8} /* (31, 25, 12) {real, imag} */,
  {32'hc2a98860, 32'h4184e68f} /* (31, 25, 11) {real, imag} */,
  {32'h40b70928, 32'h417add52} /* (31, 25, 10) {real, imag} */,
  {32'hbe045c00, 32'hc223cc4e} /* (31, 25, 9) {real, imag} */,
  {32'hc29a9203, 32'hc1b4e7b8} /* (31, 25, 8) {real, imag} */,
  {32'h424db3ea, 32'h420331d6} /* (31, 25, 7) {real, imag} */,
  {32'h3fb05340, 32'h4227d4b6} /* (31, 25, 6) {real, imag} */,
  {32'hc0de0b48, 32'hc1e48782} /* (31, 25, 5) {real, imag} */,
  {32'h425bea2d, 32'h423e147a} /* (31, 25, 4) {real, imag} */,
  {32'hc24691f8, 32'hc02508e0} /* (31, 25, 3) {real, imag} */,
  {32'hc4096ca3, 32'hc38b3aea} /* (31, 25, 2) {real, imag} */,
  {32'h4412f89d, 32'h413b7963} /* (31, 25, 1) {real, imag} */,
  {32'h43c0d8a8, 32'h00000000} /* (31, 25, 0) {real, imag} */,
  {32'h4406417a, 32'hc25612a0} /* (31, 24, 31) {real, imag} */,
  {32'hc3f531a6, 32'h436bde3f} /* (31, 24, 30) {real, imag} */,
  {32'h41306070, 32'hc2b098ee} /* (31, 24, 29) {real, imag} */,
  {32'hc1971b70, 32'hc2c4d7c7} /* (31, 24, 28) {real, imag} */,
  {32'hc2610b0b, 32'hc1df4cc0} /* (31, 24, 27) {real, imag} */,
  {32'hc22ba0bc, 32'hc28cfdb9} /* (31, 24, 26) {real, imag} */,
  {32'h420f8b63, 32'h42a1f0b6} /* (31, 24, 25) {real, imag} */,
  {32'hc30211e6, 32'h412b627e} /* (31, 24, 24) {real, imag} */,
  {32'hc239b813, 32'h42c13436} /* (31, 24, 23) {real, imag} */,
  {32'hc118cd5b, 32'hc21886a5} /* (31, 24, 22) {real, imag} */,
  {32'hc18c58d2, 32'h40e18df0} /* (31, 24, 21) {real, imag} */,
  {32'h425ba92d, 32'hc1bbbb4f} /* (31, 24, 20) {real, imag} */,
  {32'h42559846, 32'h41eaed6c} /* (31, 24, 19) {real, imag} */,
  {32'hc1de3f1b, 32'hc1ceb6a3} /* (31, 24, 18) {real, imag} */,
  {32'h4192f5dc, 32'h4266e2d3} /* (31, 24, 17) {real, imag} */,
  {32'h41e22b16, 32'h00000000} /* (31, 24, 16) {real, imag} */,
  {32'h4192f5dc, 32'hc266e2d3} /* (31, 24, 15) {real, imag} */,
  {32'hc1de3f1b, 32'h41ceb6a3} /* (31, 24, 14) {real, imag} */,
  {32'h42559846, 32'hc1eaed6c} /* (31, 24, 13) {real, imag} */,
  {32'h425ba92d, 32'h41bbbb4f} /* (31, 24, 12) {real, imag} */,
  {32'hc18c58d2, 32'hc0e18df0} /* (31, 24, 11) {real, imag} */,
  {32'hc118cd5b, 32'h421886a5} /* (31, 24, 10) {real, imag} */,
  {32'hc239b813, 32'hc2c13436} /* (31, 24, 9) {real, imag} */,
  {32'hc30211e6, 32'hc12b627e} /* (31, 24, 8) {real, imag} */,
  {32'h420f8b63, 32'hc2a1f0b6} /* (31, 24, 7) {real, imag} */,
  {32'hc22ba0bc, 32'h428cfdb9} /* (31, 24, 6) {real, imag} */,
  {32'hc2610b0b, 32'h41df4cc0} /* (31, 24, 5) {real, imag} */,
  {32'hc1971b70, 32'h42c4d7c7} /* (31, 24, 4) {real, imag} */,
  {32'h41306070, 32'h42b098ee} /* (31, 24, 3) {real, imag} */,
  {32'hc3f531a6, 32'hc36bde3f} /* (31, 24, 2) {real, imag} */,
  {32'h4406417a, 32'h425612a0} /* (31, 24, 1) {real, imag} */,
  {32'h4410df63, 32'h00000000} /* (31, 24, 0) {real, imag} */,
  {32'h43f647d1, 32'hc13006bd} /* (31, 23, 31) {real, imag} */,
  {32'hc3b673b1, 32'h433991ae} /* (31, 23, 30) {real, imag} */,
  {32'h43068e10, 32'h402c2780} /* (31, 23, 29) {real, imag} */,
  {32'hc1bb6e2a, 32'hc1fa569e} /* (31, 23, 28) {real, imag} */,
  {32'hc2d53cb8, 32'h41c0f2ba} /* (31, 23, 27) {real, imag} */,
  {32'hc23e7b46, 32'h428585ba} /* (31, 23, 26) {real, imag} */,
  {32'hc25b0809, 32'hc2553b1e} /* (31, 23, 25) {real, imag} */,
  {32'hc28ac656, 32'h42169bda} /* (31, 23, 24) {real, imag} */,
  {32'hc240f13b, 32'h4140f607} /* (31, 23, 23) {real, imag} */,
  {32'h42b73b90, 32'h42072ef4} /* (31, 23, 22) {real, imag} */,
  {32'h42849aec, 32'h4207450f} /* (31, 23, 21) {real, imag} */,
  {32'hc1f3fde6, 32'h41aa1068} /* (31, 23, 20) {real, imag} */,
  {32'h3f9e3540, 32'h421f063d} /* (31, 23, 19) {real, imag} */,
  {32'h420ab34a, 32'h4167aa24} /* (31, 23, 18) {real, imag} */,
  {32'h42534148, 32'h41c406f2} /* (31, 23, 17) {real, imag} */,
  {32'hc1a5f832, 32'h00000000} /* (31, 23, 16) {real, imag} */,
  {32'h42534148, 32'hc1c406f2} /* (31, 23, 15) {real, imag} */,
  {32'h420ab34a, 32'hc167aa24} /* (31, 23, 14) {real, imag} */,
  {32'h3f9e3540, 32'hc21f063d} /* (31, 23, 13) {real, imag} */,
  {32'hc1f3fde6, 32'hc1aa1068} /* (31, 23, 12) {real, imag} */,
  {32'h42849aec, 32'hc207450f} /* (31, 23, 11) {real, imag} */,
  {32'h42b73b90, 32'hc2072ef4} /* (31, 23, 10) {real, imag} */,
  {32'hc240f13b, 32'hc140f607} /* (31, 23, 9) {real, imag} */,
  {32'hc28ac656, 32'hc2169bda} /* (31, 23, 8) {real, imag} */,
  {32'hc25b0809, 32'h42553b1e} /* (31, 23, 7) {real, imag} */,
  {32'hc23e7b46, 32'hc28585ba} /* (31, 23, 6) {real, imag} */,
  {32'hc2d53cb8, 32'hc1c0f2ba} /* (31, 23, 5) {real, imag} */,
  {32'hc1bb6e2a, 32'h41fa569e} /* (31, 23, 4) {real, imag} */,
  {32'h43068e10, 32'hc02c2780} /* (31, 23, 3) {real, imag} */,
  {32'hc3b673b1, 32'hc33991ae} /* (31, 23, 2) {real, imag} */,
  {32'h43f647d1, 32'h413006bd} /* (31, 23, 1) {real, imag} */,
  {32'h4420dac0, 32'h00000000} /* (31, 23, 0) {real, imag} */,
  {32'h43a6460f, 32'h42f438b6} /* (31, 22, 31) {real, imag} */,
  {32'hc3b334dc, 32'h4380e432} /* (31, 22, 30) {real, imag} */,
  {32'h4368f4ce, 32'h4318044d} /* (31, 22, 29) {real, imag} */,
  {32'h420aad9a, 32'hc2028878} /* (31, 22, 28) {real, imag} */,
  {32'hc31b7fba, 32'h425bd2de} /* (31, 22, 27) {real, imag} */,
  {32'hc287e79c, 32'h41f0307b} /* (31, 22, 26) {real, imag} */,
  {32'h42a434da, 32'hc296c9c0} /* (31, 22, 25) {real, imag} */,
  {32'hc26c099f, 32'h4257184d} /* (31, 22, 24) {real, imag} */,
  {32'h3fc49490, 32'h41c88ded} /* (31, 22, 23) {real, imag} */,
  {32'hc1d13d1c, 32'h3f8f26d0} /* (31, 22, 22) {real, imag} */,
  {32'h4213e204, 32'h419bacec} /* (31, 22, 21) {real, imag} */,
  {32'hc290c03f, 32'hc159bbaf} /* (31, 22, 20) {real, imag} */,
  {32'h4243ed7c, 32'h40b8d0d8} /* (31, 22, 19) {real, imag} */,
  {32'h42321282, 32'hc29f0994} /* (31, 22, 18) {real, imag} */,
  {32'h427cb2c3, 32'hc1978318} /* (31, 22, 17) {real, imag} */,
  {32'h423e859c, 32'h00000000} /* (31, 22, 16) {real, imag} */,
  {32'h427cb2c3, 32'h41978318} /* (31, 22, 15) {real, imag} */,
  {32'h42321282, 32'h429f0994} /* (31, 22, 14) {real, imag} */,
  {32'h4243ed7c, 32'hc0b8d0d8} /* (31, 22, 13) {real, imag} */,
  {32'hc290c03f, 32'h4159bbaf} /* (31, 22, 12) {real, imag} */,
  {32'h4213e204, 32'hc19bacec} /* (31, 22, 11) {real, imag} */,
  {32'hc1d13d1c, 32'hbf8f26d0} /* (31, 22, 10) {real, imag} */,
  {32'h3fc49490, 32'hc1c88ded} /* (31, 22, 9) {real, imag} */,
  {32'hc26c099f, 32'hc257184d} /* (31, 22, 8) {real, imag} */,
  {32'h42a434da, 32'h4296c9c0} /* (31, 22, 7) {real, imag} */,
  {32'hc287e79c, 32'hc1f0307b} /* (31, 22, 6) {real, imag} */,
  {32'hc31b7fba, 32'hc25bd2de} /* (31, 22, 5) {real, imag} */,
  {32'h420aad9a, 32'h42028878} /* (31, 22, 4) {real, imag} */,
  {32'h4368f4ce, 32'hc318044d} /* (31, 22, 3) {real, imag} */,
  {32'hc3b334dc, 32'hc380e432} /* (31, 22, 2) {real, imag} */,
  {32'h43a6460f, 32'hc2f438b6} /* (31, 22, 1) {real, imag} */,
  {32'h43ed0004, 32'h00000000} /* (31, 22, 0) {real, imag} */,
  {32'h40064600, 32'h42cd1da6} /* (31, 21, 31) {real, imag} */,
  {32'hc3250786, 32'h42154c93} /* (31, 21, 30) {real, imag} */,
  {32'h42dd6a28, 32'h42910ff2} /* (31, 21, 29) {real, imag} */,
  {32'hc2b55600, 32'hc26c0395} /* (31, 21, 28) {real, imag} */,
  {32'hc29781f8, 32'hc04055c8} /* (31, 21, 27) {real, imag} */,
  {32'hc26d730e, 32'hc1837aa3} /* (31, 21, 26) {real, imag} */,
  {32'hc1f02309, 32'h41f5f784} /* (31, 21, 25) {real, imag} */,
  {32'h421a849a, 32'hc166216c} /* (31, 21, 24) {real, imag} */,
  {32'hc2a657f4, 32'h4223c0ad} /* (31, 21, 23) {real, imag} */,
  {32'h417eadc3, 32'hc212f304} /* (31, 21, 22) {real, imag} */,
  {32'h40e91dc8, 32'h420db374} /* (31, 21, 21) {real, imag} */,
  {32'hc246b9ae, 32'hc0bd1b9c} /* (31, 21, 20) {real, imag} */,
  {32'hc2895178, 32'h42324d58} /* (31, 21, 19) {real, imag} */,
  {32'h40c65ec8, 32'h41813829} /* (31, 21, 18) {real, imag} */,
  {32'h41a57d30, 32'hc15a6966} /* (31, 21, 17) {real, imag} */,
  {32'h41f369b1, 32'h00000000} /* (31, 21, 16) {real, imag} */,
  {32'h41a57d30, 32'h415a6966} /* (31, 21, 15) {real, imag} */,
  {32'h40c65ec8, 32'hc1813829} /* (31, 21, 14) {real, imag} */,
  {32'hc2895178, 32'hc2324d58} /* (31, 21, 13) {real, imag} */,
  {32'hc246b9ae, 32'h40bd1b9c} /* (31, 21, 12) {real, imag} */,
  {32'h40e91dc8, 32'hc20db374} /* (31, 21, 11) {real, imag} */,
  {32'h417eadc3, 32'h4212f304} /* (31, 21, 10) {real, imag} */,
  {32'hc2a657f4, 32'hc223c0ad} /* (31, 21, 9) {real, imag} */,
  {32'h421a849a, 32'h4166216c} /* (31, 21, 8) {real, imag} */,
  {32'hc1f02309, 32'hc1f5f784} /* (31, 21, 7) {real, imag} */,
  {32'hc26d730e, 32'h41837aa3} /* (31, 21, 6) {real, imag} */,
  {32'hc29781f8, 32'h404055c8} /* (31, 21, 5) {real, imag} */,
  {32'hc2b55600, 32'h426c0395} /* (31, 21, 4) {real, imag} */,
  {32'h42dd6a28, 32'hc2910ff2} /* (31, 21, 3) {real, imag} */,
  {32'hc3250786, 32'hc2154c93} /* (31, 21, 2) {real, imag} */,
  {32'h40064600, 32'hc2cd1da6} /* (31, 21, 1) {real, imag} */,
  {32'h4329b110, 32'h00000000} /* (31, 21, 0) {real, imag} */,
  {32'hc3f7b100, 32'h428307fe} /* (31, 20, 31) {real, imag} */,
  {32'h432fa0e0, 32'hc34c94ec} /* (31, 20, 30) {real, imag} */,
  {32'h42a985e1, 32'h42bb88da} /* (31, 20, 29) {real, imag} */,
  {32'hc330be2d, 32'h422f58c5} /* (31, 20, 28) {real, imag} */,
  {32'h42828483, 32'h4121c40c} /* (31, 20, 27) {real, imag} */,
  {32'hbdea77c0, 32'hc2a2feb8} /* (31, 20, 26) {real, imag} */,
  {32'h420babc8, 32'hc22b65bf} /* (31, 20, 25) {real, imag} */,
  {32'h3fdb53c0, 32'h421ea775} /* (31, 20, 24) {real, imag} */,
  {32'hc21212b6, 32'h42354348} /* (31, 20, 23) {real, imag} */,
  {32'h41b4fc42, 32'hc2695d8c} /* (31, 20, 22) {real, imag} */,
  {32'hc29a3e4e, 32'hc24e9ebd} /* (31, 20, 21) {real, imag} */,
  {32'hc29eedac, 32'hc15690e8} /* (31, 20, 20) {real, imag} */,
  {32'h41dceefe, 32'h429ed2e1} /* (31, 20, 19) {real, imag} */,
  {32'hc10bb260, 32'hc0f44d30} /* (31, 20, 18) {real, imag} */,
  {32'hbeee0c80, 32'h424f0855} /* (31, 20, 17) {real, imag} */,
  {32'hc19f84a7, 32'h00000000} /* (31, 20, 16) {real, imag} */,
  {32'hbeee0c80, 32'hc24f0855} /* (31, 20, 15) {real, imag} */,
  {32'hc10bb260, 32'h40f44d30} /* (31, 20, 14) {real, imag} */,
  {32'h41dceefe, 32'hc29ed2e1} /* (31, 20, 13) {real, imag} */,
  {32'hc29eedac, 32'h415690e8} /* (31, 20, 12) {real, imag} */,
  {32'hc29a3e4e, 32'h424e9ebd} /* (31, 20, 11) {real, imag} */,
  {32'h41b4fc42, 32'h42695d8c} /* (31, 20, 10) {real, imag} */,
  {32'hc21212b6, 32'hc2354348} /* (31, 20, 9) {real, imag} */,
  {32'h3fdb53c0, 32'hc21ea775} /* (31, 20, 8) {real, imag} */,
  {32'h420babc8, 32'h422b65bf} /* (31, 20, 7) {real, imag} */,
  {32'hbdea77c0, 32'h42a2feb8} /* (31, 20, 6) {real, imag} */,
  {32'h42828483, 32'hc121c40c} /* (31, 20, 5) {real, imag} */,
  {32'hc330be2d, 32'hc22f58c5} /* (31, 20, 4) {real, imag} */,
  {32'h42a985e1, 32'hc2bb88da} /* (31, 20, 3) {real, imag} */,
  {32'h432fa0e0, 32'h434c94ec} /* (31, 20, 2) {real, imag} */,
  {32'hc3f7b100, 32'hc28307fe} /* (31, 20, 1) {real, imag} */,
  {32'hc3ae5500, 32'h00000000} /* (31, 20, 0) {real, imag} */,
  {32'hc44afe9a, 32'h421efef0} /* (31, 19, 31) {real, imag} */,
  {32'h43b303e8, 32'hc337f0c8} /* (31, 19, 30) {real, imag} */,
  {32'hc12c4bc6, 32'h428c467a} /* (31, 19, 29) {real, imag} */,
  {32'hc33e77db, 32'hc285d5ee} /* (31, 19, 28) {real, imag} */,
  {32'h42cdb140, 32'hc2dbd229} /* (31, 19, 27) {real, imag} */,
  {32'h41848964, 32'h426ad2b9} /* (31, 19, 26) {real, imag} */,
  {32'hc194d3ae, 32'h42766f9c} /* (31, 19, 25) {real, imag} */,
  {32'hc235f6ba, 32'hc1b36c10} /* (31, 19, 24) {real, imag} */,
  {32'h41080985, 32'h41fcc8b0} /* (31, 19, 23) {real, imag} */,
  {32'hc25c9120, 32'hc2966fc4} /* (31, 19, 22) {real, imag} */,
  {32'hc25cd2f1, 32'h41dc6ec1} /* (31, 19, 21) {real, imag} */,
  {32'h4216d3dc, 32'hc2af4f3d} /* (31, 19, 20) {real, imag} */,
  {32'hc1df72ca, 32'hc2931579} /* (31, 19, 19) {real, imag} */,
  {32'hc18781bb, 32'hc2d922b2} /* (31, 19, 18) {real, imag} */,
  {32'hc0a33488, 32'h41efc944} /* (31, 19, 17) {real, imag} */,
  {32'h41bfe1d6, 32'h00000000} /* (31, 19, 16) {real, imag} */,
  {32'hc0a33488, 32'hc1efc944} /* (31, 19, 15) {real, imag} */,
  {32'hc18781bb, 32'h42d922b2} /* (31, 19, 14) {real, imag} */,
  {32'hc1df72ca, 32'h42931579} /* (31, 19, 13) {real, imag} */,
  {32'h4216d3dc, 32'h42af4f3d} /* (31, 19, 12) {real, imag} */,
  {32'hc25cd2f1, 32'hc1dc6ec1} /* (31, 19, 11) {real, imag} */,
  {32'hc25c9120, 32'h42966fc4} /* (31, 19, 10) {real, imag} */,
  {32'h41080985, 32'hc1fcc8b0} /* (31, 19, 9) {real, imag} */,
  {32'hc235f6ba, 32'h41b36c10} /* (31, 19, 8) {real, imag} */,
  {32'hc194d3ae, 32'hc2766f9c} /* (31, 19, 7) {real, imag} */,
  {32'h41848964, 32'hc26ad2b9} /* (31, 19, 6) {real, imag} */,
  {32'h42cdb140, 32'h42dbd229} /* (31, 19, 5) {real, imag} */,
  {32'hc33e77db, 32'h4285d5ee} /* (31, 19, 4) {real, imag} */,
  {32'hc12c4bc6, 32'hc28c467a} /* (31, 19, 3) {real, imag} */,
  {32'h43b303e8, 32'h4337f0c8} /* (31, 19, 2) {real, imag} */,
  {32'hc44afe9a, 32'hc21efef0} /* (31, 19, 1) {real, imag} */,
  {32'hc3eed135, 32'h00000000} /* (31, 19, 0) {real, imag} */,
  {32'hc453a90a, 32'hc22d3beb} /* (31, 18, 31) {real, imag} */,
  {32'h43a03c6c, 32'hc306c17a} /* (31, 18, 30) {real, imag} */,
  {32'hc22b3bb6, 32'h42bd2c4d} /* (31, 18, 29) {real, imag} */,
  {32'hc38776ff, 32'h41e9a8d5} /* (31, 18, 28) {real, imag} */,
  {32'h43048b1f, 32'hc261865e} /* (31, 18, 27) {real, imag} */,
  {32'h40a99dec, 32'hc0011e40} /* (31, 18, 26) {real, imag} */,
  {32'h41778805, 32'hc12edf16} /* (31, 18, 25) {real, imag} */,
  {32'h424f3ce0, 32'h41064c1c} /* (31, 18, 24) {real, imag} */,
  {32'h400b9bb8, 32'h4244e70c} /* (31, 18, 23) {real, imag} */,
  {32'h420a8487, 32'hc1c0de60} /* (31, 18, 22) {real, imag} */,
  {32'h40e7ecac, 32'h419678f2} /* (31, 18, 21) {real, imag} */,
  {32'h426824eb, 32'h4163dc8c} /* (31, 18, 20) {real, imag} */,
  {32'h42bf60cd, 32'h41122e40} /* (31, 18, 19) {real, imag} */,
  {32'hc0872e22, 32'hc14bacfe} /* (31, 18, 18) {real, imag} */,
  {32'h41328088, 32'h41bcda76} /* (31, 18, 17) {real, imag} */,
  {32'h414313fb, 32'h00000000} /* (31, 18, 16) {real, imag} */,
  {32'h41328088, 32'hc1bcda76} /* (31, 18, 15) {real, imag} */,
  {32'hc0872e22, 32'h414bacfe} /* (31, 18, 14) {real, imag} */,
  {32'h42bf60cd, 32'hc1122e40} /* (31, 18, 13) {real, imag} */,
  {32'h426824eb, 32'hc163dc8c} /* (31, 18, 12) {real, imag} */,
  {32'h40e7ecac, 32'hc19678f2} /* (31, 18, 11) {real, imag} */,
  {32'h420a8487, 32'h41c0de60} /* (31, 18, 10) {real, imag} */,
  {32'h400b9bb8, 32'hc244e70c} /* (31, 18, 9) {real, imag} */,
  {32'h424f3ce0, 32'hc1064c1c} /* (31, 18, 8) {real, imag} */,
  {32'h41778805, 32'h412edf16} /* (31, 18, 7) {real, imag} */,
  {32'h40a99dec, 32'h40011e40} /* (31, 18, 6) {real, imag} */,
  {32'h43048b1f, 32'h4261865e} /* (31, 18, 5) {real, imag} */,
  {32'hc38776ff, 32'hc1e9a8d5} /* (31, 18, 4) {real, imag} */,
  {32'hc22b3bb6, 32'hc2bd2c4d} /* (31, 18, 3) {real, imag} */,
  {32'h43a03c6c, 32'h4306c17a} /* (31, 18, 2) {real, imag} */,
  {32'hc453a90a, 32'h422d3beb} /* (31, 18, 1) {real, imag} */,
  {32'hc3b518bb, 32'h00000000} /* (31, 18, 0) {real, imag} */,
  {32'hc4532f85, 32'hc3176cf1} /* (31, 17, 31) {real, imag} */,
  {32'h4381587c, 32'hc27b08a0} /* (31, 17, 30) {real, imag} */,
  {32'hc269a700, 32'h40e46aa8} /* (31, 17, 29) {real, imag} */,
  {32'hc3186532, 32'h3fb82828} /* (31, 17, 28) {real, imag} */,
  {32'h42ce08bb, 32'hc23733fb} /* (31, 17, 27) {real, imag} */,
  {32'hc136faf3, 32'hc208cd2b} /* (31, 17, 26) {real, imag} */,
  {32'hc2722c02, 32'h426200cd} /* (31, 17, 25) {real, imag} */,
  {32'h41e6f0c0, 32'hc2929768} /* (31, 17, 24) {real, imag} */,
  {32'h41268e9e, 32'hc2462382} /* (31, 17, 23) {real, imag} */,
  {32'hc1bf4967, 32'h4201ca11} /* (31, 17, 22) {real, imag} */,
  {32'h4271d9ce, 32'hc233d88f} /* (31, 17, 21) {real, imag} */,
  {32'hc28fe250, 32'hc1745ab7} /* (31, 17, 20) {real, imag} */,
  {32'h41df2d32, 32'h4082b338} /* (31, 17, 19) {real, imag} */,
  {32'h421d2ba2, 32'hc271fb9d} /* (31, 17, 18) {real, imag} */,
  {32'h40edc480, 32'h40829f34} /* (31, 17, 17) {real, imag} */,
  {32'h4258e79f, 32'h00000000} /* (31, 17, 16) {real, imag} */,
  {32'h40edc480, 32'hc0829f34} /* (31, 17, 15) {real, imag} */,
  {32'h421d2ba2, 32'h4271fb9d} /* (31, 17, 14) {real, imag} */,
  {32'h41df2d32, 32'hc082b338} /* (31, 17, 13) {real, imag} */,
  {32'hc28fe250, 32'h41745ab7} /* (31, 17, 12) {real, imag} */,
  {32'h4271d9ce, 32'h4233d88f} /* (31, 17, 11) {real, imag} */,
  {32'hc1bf4967, 32'hc201ca11} /* (31, 17, 10) {real, imag} */,
  {32'h41268e9e, 32'h42462382} /* (31, 17, 9) {real, imag} */,
  {32'h41e6f0c0, 32'h42929768} /* (31, 17, 8) {real, imag} */,
  {32'hc2722c02, 32'hc26200cd} /* (31, 17, 7) {real, imag} */,
  {32'hc136faf3, 32'h4208cd2b} /* (31, 17, 6) {real, imag} */,
  {32'h42ce08bb, 32'h423733fb} /* (31, 17, 5) {real, imag} */,
  {32'hc3186532, 32'hbfb82828} /* (31, 17, 4) {real, imag} */,
  {32'hc269a700, 32'hc0e46aa8} /* (31, 17, 3) {real, imag} */,
  {32'h4381587c, 32'h427b08a0} /* (31, 17, 2) {real, imag} */,
  {32'hc4532f85, 32'h43176cf1} /* (31, 17, 1) {real, imag} */,
  {32'hc3bf0c9a, 32'h00000000} /* (31, 17, 0) {real, imag} */,
  {32'hc442bdd8, 32'hc326ac52} /* (31, 16, 31) {real, imag} */,
  {32'h43a17533, 32'hc2e7971e} /* (31, 16, 30) {real, imag} */,
  {32'hc2603081, 32'h428cd869} /* (31, 16, 29) {real, imag} */,
  {32'hc30bbbb5, 32'h40bbe650} /* (31, 16, 28) {real, imag} */,
  {32'h42d03b02, 32'h40c2f800} /* (31, 16, 27) {real, imag} */,
  {32'hc233c628, 32'h41c79be1} /* (31, 16, 26) {real, imag} */,
  {32'hc26106e4, 32'hc2763793} /* (31, 16, 25) {real, imag} */,
  {32'h42c069ba, 32'hc281eae8} /* (31, 16, 24) {real, imag} */,
  {32'hc20885d4, 32'hc21be1f0} /* (31, 16, 23) {real, imag} */,
  {32'hc1a074f4, 32'h400d7f68} /* (31, 16, 22) {real, imag} */,
  {32'hc1b54d5a, 32'hc14e14f7} /* (31, 16, 21) {real, imag} */,
  {32'hc2223446, 32'hc22652b5} /* (31, 16, 20) {real, imag} */,
  {32'h41d8baf6, 32'hc1a1def6} /* (31, 16, 19) {real, imag} */,
  {32'h41393810, 32'h41f9e8f6} /* (31, 16, 18) {real, imag} */,
  {32'hc22b38ab, 32'h41844c1e} /* (31, 16, 17) {real, imag} */,
  {32'h4203f96d, 32'h00000000} /* (31, 16, 16) {real, imag} */,
  {32'hc22b38ab, 32'hc1844c1e} /* (31, 16, 15) {real, imag} */,
  {32'h41393810, 32'hc1f9e8f6} /* (31, 16, 14) {real, imag} */,
  {32'h41d8baf6, 32'h41a1def6} /* (31, 16, 13) {real, imag} */,
  {32'hc2223446, 32'h422652b5} /* (31, 16, 12) {real, imag} */,
  {32'hc1b54d5a, 32'h414e14f7} /* (31, 16, 11) {real, imag} */,
  {32'hc1a074f4, 32'hc00d7f68} /* (31, 16, 10) {real, imag} */,
  {32'hc20885d4, 32'h421be1f0} /* (31, 16, 9) {real, imag} */,
  {32'h42c069ba, 32'h4281eae8} /* (31, 16, 8) {real, imag} */,
  {32'hc26106e4, 32'h42763793} /* (31, 16, 7) {real, imag} */,
  {32'hc233c628, 32'hc1c79be1} /* (31, 16, 6) {real, imag} */,
  {32'h42d03b02, 32'hc0c2f800} /* (31, 16, 5) {real, imag} */,
  {32'hc30bbbb5, 32'hc0bbe650} /* (31, 16, 4) {real, imag} */,
  {32'hc2603081, 32'hc28cd869} /* (31, 16, 3) {real, imag} */,
  {32'h43a17533, 32'h42e7971e} /* (31, 16, 2) {real, imag} */,
  {32'hc442bdd8, 32'h4326ac52} /* (31, 16, 1) {real, imag} */,
  {32'hc4023467, 32'h00000000} /* (31, 16, 0) {real, imag} */,
  {32'hc42bbffb, 32'hc30edc53} /* (31, 15, 31) {real, imag} */,
  {32'h4391341c, 32'hc2d51164} /* (31, 15, 30) {real, imag} */,
  {32'hc26c305c, 32'h42b07aac} /* (31, 15, 29) {real, imag} */,
  {32'hc28e9a53, 32'h41862a0e} /* (31, 15, 28) {real, imag} */,
  {32'h42d8dff9, 32'h4290fc28} /* (31, 15, 27) {real, imag} */,
  {32'h3ea1db20, 32'hc137dce0} /* (31, 15, 26) {real, imag} */,
  {32'h4100f470, 32'hc2061df9} /* (31, 15, 25) {real, imag} */,
  {32'h41e4dc04, 32'hc196bb5e} /* (31, 15, 24) {real, imag} */,
  {32'h41e949a1, 32'h419433b8} /* (31, 15, 23) {real, imag} */,
  {32'hc18a4931, 32'hc29fd9d6} /* (31, 15, 22) {real, imag} */,
  {32'h405c40e0, 32'hc1f359f6} /* (31, 15, 21) {real, imag} */,
  {32'h42a158a0, 32'h4195425a} /* (31, 15, 20) {real, imag} */,
  {32'h427f82cd, 32'h423697c1} /* (31, 15, 19) {real, imag} */,
  {32'h4168b04b, 32'h41a889d6} /* (31, 15, 18) {real, imag} */,
  {32'h4227d79a, 32'h420f53ae} /* (31, 15, 17) {real, imag} */,
  {32'h41eee59a, 32'h00000000} /* (31, 15, 16) {real, imag} */,
  {32'h4227d79a, 32'hc20f53ae} /* (31, 15, 15) {real, imag} */,
  {32'h4168b04b, 32'hc1a889d6} /* (31, 15, 14) {real, imag} */,
  {32'h427f82cd, 32'hc23697c1} /* (31, 15, 13) {real, imag} */,
  {32'h42a158a0, 32'hc195425a} /* (31, 15, 12) {real, imag} */,
  {32'h405c40e0, 32'h41f359f6} /* (31, 15, 11) {real, imag} */,
  {32'hc18a4931, 32'h429fd9d6} /* (31, 15, 10) {real, imag} */,
  {32'h41e949a1, 32'hc19433b8} /* (31, 15, 9) {real, imag} */,
  {32'h41e4dc04, 32'h4196bb5e} /* (31, 15, 8) {real, imag} */,
  {32'h4100f470, 32'h42061df9} /* (31, 15, 7) {real, imag} */,
  {32'h3ea1db20, 32'h4137dce0} /* (31, 15, 6) {real, imag} */,
  {32'h42d8dff9, 32'hc290fc28} /* (31, 15, 5) {real, imag} */,
  {32'hc28e9a53, 32'hc1862a0e} /* (31, 15, 4) {real, imag} */,
  {32'hc26c305c, 32'hc2b07aac} /* (31, 15, 3) {real, imag} */,
  {32'h4391341c, 32'h42d51164} /* (31, 15, 2) {real, imag} */,
  {32'hc42bbffb, 32'h430edc53} /* (31, 15, 1) {real, imag} */,
  {32'hc41853e1, 32'h00000000} /* (31, 15, 0) {real, imag} */,
  {32'hc4092f0c, 32'hc2dfca0a} /* (31, 14, 31) {real, imag} */,
  {32'h43a5ae28, 32'h419d2ad4} /* (31, 14, 30) {real, imag} */,
  {32'hc190b0a0, 32'h4229819e} /* (31, 14, 29) {real, imag} */,
  {32'h41a5f75c, 32'h426cf3f2} /* (31, 14, 28) {real, imag} */,
  {32'h42751a55, 32'h41c44e44} /* (31, 14, 27) {real, imag} */,
  {32'h421588a6, 32'hbe1b3100} /* (31, 14, 26) {real, imag} */,
  {32'hc22a3fad, 32'h4283cfb3} /* (31, 14, 25) {real, imag} */,
  {32'h4245febe, 32'hc2732423} /* (31, 14, 24) {real, imag} */,
  {32'hc0efb44c, 32'hc1787ab8} /* (31, 14, 23) {real, imag} */,
  {32'h415efb1c, 32'h41e52e08} /* (31, 14, 22) {real, imag} */,
  {32'h42829d2c, 32'h413d83c9} /* (31, 14, 21) {real, imag} */,
  {32'hc2a2105e, 32'hc0848730} /* (31, 14, 20) {real, imag} */,
  {32'hc1dfa17c, 32'hc1562d8c} /* (31, 14, 19) {real, imag} */,
  {32'hc1a598b8, 32'hc1651fb6} /* (31, 14, 18) {real, imag} */,
  {32'h40a4ac0f, 32'h41389bdc} /* (31, 14, 17) {real, imag} */,
  {32'h40cc129a, 32'h00000000} /* (31, 14, 16) {real, imag} */,
  {32'h40a4ac0f, 32'hc1389bdc} /* (31, 14, 15) {real, imag} */,
  {32'hc1a598b8, 32'h41651fb6} /* (31, 14, 14) {real, imag} */,
  {32'hc1dfa17c, 32'h41562d8c} /* (31, 14, 13) {real, imag} */,
  {32'hc2a2105e, 32'h40848730} /* (31, 14, 12) {real, imag} */,
  {32'h42829d2c, 32'hc13d83c9} /* (31, 14, 11) {real, imag} */,
  {32'h415efb1c, 32'hc1e52e08} /* (31, 14, 10) {real, imag} */,
  {32'hc0efb44c, 32'h41787ab8} /* (31, 14, 9) {real, imag} */,
  {32'h4245febe, 32'h42732423} /* (31, 14, 8) {real, imag} */,
  {32'hc22a3fad, 32'hc283cfb3} /* (31, 14, 7) {real, imag} */,
  {32'h421588a6, 32'h3e1b3100} /* (31, 14, 6) {real, imag} */,
  {32'h42751a55, 32'hc1c44e44} /* (31, 14, 5) {real, imag} */,
  {32'h41a5f75c, 32'hc26cf3f2} /* (31, 14, 4) {real, imag} */,
  {32'hc190b0a0, 32'hc229819e} /* (31, 14, 3) {real, imag} */,
  {32'h43a5ae28, 32'hc19d2ad4} /* (31, 14, 2) {real, imag} */,
  {32'hc4092f0c, 32'h42dfca0a} /* (31, 14, 1) {real, imag} */,
  {32'hc4273b1e, 32'h00000000} /* (31, 14, 0) {real, imag} */,
  {32'hc4011068, 32'hc2c48184} /* (31, 13, 31) {real, imag} */,
  {32'h43d5f904, 32'hc2b13f80} /* (31, 13, 30) {real, imag} */,
  {32'hc25bfc5e, 32'h4259dc28} /* (31, 13, 29) {real, imag} */,
  {32'hc2f03132, 32'h42026dcc} /* (31, 13, 28) {real, imag} */,
  {32'h423960db, 32'h4045e560} /* (31, 13, 27) {real, imag} */,
  {32'h4245872c, 32'hc1caf876} /* (31, 13, 26) {real, imag} */,
  {32'h420e977b, 32'h425d8dac} /* (31, 13, 25) {real, imag} */,
  {32'h416a3732, 32'hc2316052} /* (31, 13, 24) {real, imag} */,
  {32'h4101309b, 32'hc268d9fc} /* (31, 13, 23) {real, imag} */,
  {32'h42567610, 32'h41b8f926} /* (31, 13, 22) {real, imag} */,
  {32'hc0067340, 32'h4240f474} /* (31, 13, 21) {real, imag} */,
  {32'hc2932ec7, 32'hc1e69c1b} /* (31, 13, 20) {real, imag} */,
  {32'h41d7b438, 32'h4182c8bc} /* (31, 13, 19) {real, imag} */,
  {32'h3daca300, 32'h411fc4ac} /* (31, 13, 18) {real, imag} */,
  {32'h40b47050, 32'hc1a8df44} /* (31, 13, 17) {real, imag} */,
  {32'hc2345879, 32'h00000000} /* (31, 13, 16) {real, imag} */,
  {32'h40b47050, 32'h41a8df44} /* (31, 13, 15) {real, imag} */,
  {32'h3daca300, 32'hc11fc4ac} /* (31, 13, 14) {real, imag} */,
  {32'h41d7b438, 32'hc182c8bc} /* (31, 13, 13) {real, imag} */,
  {32'hc2932ec7, 32'h41e69c1b} /* (31, 13, 12) {real, imag} */,
  {32'hc0067340, 32'hc240f474} /* (31, 13, 11) {real, imag} */,
  {32'h42567610, 32'hc1b8f926} /* (31, 13, 10) {real, imag} */,
  {32'h4101309b, 32'h4268d9fc} /* (31, 13, 9) {real, imag} */,
  {32'h416a3732, 32'h42316052} /* (31, 13, 8) {real, imag} */,
  {32'h420e977b, 32'hc25d8dac} /* (31, 13, 7) {real, imag} */,
  {32'h4245872c, 32'h41caf876} /* (31, 13, 6) {real, imag} */,
  {32'h423960db, 32'hc045e560} /* (31, 13, 5) {real, imag} */,
  {32'hc2f03132, 32'hc2026dcc} /* (31, 13, 4) {real, imag} */,
  {32'hc25bfc5e, 32'hc259dc28} /* (31, 13, 3) {real, imag} */,
  {32'h43d5f904, 32'h42b13f80} /* (31, 13, 2) {real, imag} */,
  {32'hc4011068, 32'h42c48184} /* (31, 13, 1) {real, imag} */,
  {32'hc430a0d8, 32'h00000000} /* (31, 13, 0) {real, imag} */,
  {32'hc3f64d92, 32'hbd3e3000} /* (31, 12, 31) {real, imag} */,
  {32'h43c075d0, 32'hc2938c41} /* (31, 12, 30) {real, imag} */,
  {32'hc291c6b3, 32'h428c2a42} /* (31, 12, 29) {real, imag} */,
  {32'hc2dece3e, 32'h414cc33d} /* (31, 12, 28) {real, imag} */,
  {32'h3fb21b30, 32'hc2ba70e4} /* (31, 12, 27) {real, imag} */,
  {32'hbf7ef8c8, 32'h4176bc74} /* (31, 12, 26) {real, imag} */,
  {32'hc2c6af64, 32'h4284b6c8} /* (31, 12, 25) {real, imag} */,
  {32'h42b2f17f, 32'hc0bad4c8} /* (31, 12, 24) {real, imag} */,
  {32'h422bdd5e, 32'hc26dda90} /* (31, 12, 23) {real, imag} */,
  {32'h40efadca, 32'hc2370a74} /* (31, 12, 22) {real, imag} */,
  {32'hc258fb71, 32'hc1b72c56} /* (31, 12, 21) {real, imag} */,
  {32'h3fb375a0, 32'hc062bd22} /* (31, 12, 20) {real, imag} */,
  {32'h41260ae4, 32'hc2a32895} /* (31, 12, 19) {real, imag} */,
  {32'h42db4424, 32'hc16ceb10} /* (31, 12, 18) {real, imag} */,
  {32'hc2158ed2, 32'hc188f942} /* (31, 12, 17) {real, imag} */,
  {32'hc231a466, 32'h00000000} /* (31, 12, 16) {real, imag} */,
  {32'hc2158ed2, 32'h4188f942} /* (31, 12, 15) {real, imag} */,
  {32'h42db4424, 32'h416ceb10} /* (31, 12, 14) {real, imag} */,
  {32'h41260ae4, 32'h42a32895} /* (31, 12, 13) {real, imag} */,
  {32'h3fb375a0, 32'h4062bd22} /* (31, 12, 12) {real, imag} */,
  {32'hc258fb71, 32'h41b72c56} /* (31, 12, 11) {real, imag} */,
  {32'h40efadca, 32'h42370a74} /* (31, 12, 10) {real, imag} */,
  {32'h422bdd5e, 32'h426dda90} /* (31, 12, 9) {real, imag} */,
  {32'h42b2f17f, 32'h40bad4c8} /* (31, 12, 8) {real, imag} */,
  {32'hc2c6af64, 32'hc284b6c8} /* (31, 12, 7) {real, imag} */,
  {32'hbf7ef8c8, 32'hc176bc74} /* (31, 12, 6) {real, imag} */,
  {32'h3fb21b30, 32'h42ba70e4} /* (31, 12, 5) {real, imag} */,
  {32'hc2dece3e, 32'hc14cc33d} /* (31, 12, 4) {real, imag} */,
  {32'hc291c6b3, 32'hc28c2a42} /* (31, 12, 3) {real, imag} */,
  {32'h43c075d0, 32'h42938c41} /* (31, 12, 2) {real, imag} */,
  {32'hc3f64d92, 32'h3d3e3000} /* (31, 12, 1) {real, imag} */,
  {32'hc428df90, 32'h00000000} /* (31, 12, 0) {real, imag} */,
  {32'hc382e638, 32'h41a48a98} /* (31, 11, 31) {real, imag} */,
  {32'h4378da9a, 32'h420c08a1} /* (31, 11, 30) {real, imag} */,
  {32'hc2458fed, 32'hc1a91446} /* (31, 11, 29) {real, imag} */,
  {32'h4209f048, 32'h42763eff} /* (31, 11, 28) {real, imag} */,
  {32'h42b8a14e, 32'hc285574c} /* (31, 11, 27) {real, imag} */,
  {32'h4104209a, 32'h4251ccd4} /* (31, 11, 26) {real, imag} */,
  {32'hc290824f, 32'hbffeb220} /* (31, 11, 25) {real, imag} */,
  {32'h4273202a, 32'h411ad730} /* (31, 11, 24) {real, imag} */,
  {32'h428f3cd2, 32'hc2085fcf} /* (31, 11, 23) {real, imag} */,
  {32'h41a27fdc, 32'h426118b4} /* (31, 11, 22) {real, imag} */,
  {32'h42c7f3e0, 32'hc25f9cee} /* (31, 11, 21) {real, imag} */,
  {32'hc2bf5ac1, 32'h4210df72} /* (31, 11, 20) {real, imag} */,
  {32'hc28192cc, 32'hc2255c5a} /* (31, 11, 19) {real, imag} */,
  {32'hc1a7cb2a, 32'h40319e58} /* (31, 11, 18) {real, imag} */,
  {32'hc02ec194, 32'hc1adca19} /* (31, 11, 17) {real, imag} */,
  {32'h421ffa9c, 32'h00000000} /* (31, 11, 16) {real, imag} */,
  {32'hc02ec194, 32'h41adca19} /* (31, 11, 15) {real, imag} */,
  {32'hc1a7cb2a, 32'hc0319e58} /* (31, 11, 14) {real, imag} */,
  {32'hc28192cc, 32'h42255c5a} /* (31, 11, 13) {real, imag} */,
  {32'hc2bf5ac1, 32'hc210df72} /* (31, 11, 12) {real, imag} */,
  {32'h42c7f3e0, 32'h425f9cee} /* (31, 11, 11) {real, imag} */,
  {32'h41a27fdc, 32'hc26118b4} /* (31, 11, 10) {real, imag} */,
  {32'h428f3cd2, 32'h42085fcf} /* (31, 11, 9) {real, imag} */,
  {32'h4273202a, 32'hc11ad730} /* (31, 11, 8) {real, imag} */,
  {32'hc290824f, 32'h3ffeb220} /* (31, 11, 7) {real, imag} */,
  {32'h4104209a, 32'hc251ccd4} /* (31, 11, 6) {real, imag} */,
  {32'h42b8a14e, 32'h4285574c} /* (31, 11, 5) {real, imag} */,
  {32'h4209f048, 32'hc2763eff} /* (31, 11, 4) {real, imag} */,
  {32'hc2458fed, 32'h41a91446} /* (31, 11, 3) {real, imag} */,
  {32'h4378da9a, 32'hc20c08a1} /* (31, 11, 2) {real, imag} */,
  {32'hc382e638, 32'hc1a48a98} /* (31, 11, 1) {real, imag} */,
  {32'hc3a1e3c1, 32'h00000000} /* (31, 11, 0) {real, imag} */,
  {32'h439c28bd, 32'h423513fb} /* (31, 10, 31) {real, imag} */,
  {32'hc327fb8b, 32'h42ec3bea} /* (31, 10, 30) {real, imag} */,
  {32'h424685e8, 32'hc2eeecde} /* (31, 10, 29) {real, imag} */,
  {32'h42ac3c32, 32'h41b8537f} /* (31, 10, 28) {real, imag} */,
  {32'h409a9b50, 32'hc30d3a9e} /* (31, 10, 27) {real, imag} */,
  {32'hc18f6dba, 32'h41e77efb} /* (31, 10, 26) {real, imag} */,
  {32'hc1f75c40, 32'hc2d95afc} /* (31, 10, 25) {real, imag} */,
  {32'h4130bcd4, 32'h4250cfd3} /* (31, 10, 24) {real, imag} */,
  {32'hc272a842, 32'hc272887e} /* (31, 10, 23) {real, imag} */,
  {32'hc24f351a, 32'h42527988} /* (31, 10, 22) {real, imag} */,
  {32'hc2636dc8, 32'hc29f035d} /* (31, 10, 21) {real, imag} */,
  {32'hc220d244, 32'h4151dabb} /* (31, 10, 20) {real, imag} */,
  {32'hc29660ec, 32'hc0a17be8} /* (31, 10, 19) {real, imag} */,
  {32'h4301fe72, 32'h423861e5} /* (31, 10, 18) {real, imag} */,
  {32'hc23d46e3, 32'hc25ee7de} /* (31, 10, 17) {real, imag} */,
  {32'h40e9d420, 32'h00000000} /* (31, 10, 16) {real, imag} */,
  {32'hc23d46e3, 32'h425ee7de} /* (31, 10, 15) {real, imag} */,
  {32'h4301fe72, 32'hc23861e5} /* (31, 10, 14) {real, imag} */,
  {32'hc29660ec, 32'h40a17be8} /* (31, 10, 13) {real, imag} */,
  {32'hc220d244, 32'hc151dabb} /* (31, 10, 12) {real, imag} */,
  {32'hc2636dc8, 32'h429f035d} /* (31, 10, 11) {real, imag} */,
  {32'hc24f351a, 32'hc2527988} /* (31, 10, 10) {real, imag} */,
  {32'hc272a842, 32'h4272887e} /* (31, 10, 9) {real, imag} */,
  {32'h4130bcd4, 32'hc250cfd3} /* (31, 10, 8) {real, imag} */,
  {32'hc1f75c40, 32'h42d95afc} /* (31, 10, 7) {real, imag} */,
  {32'hc18f6dba, 32'hc1e77efb} /* (31, 10, 6) {real, imag} */,
  {32'h409a9b50, 32'h430d3a9e} /* (31, 10, 5) {real, imag} */,
  {32'h42ac3c32, 32'hc1b8537f} /* (31, 10, 4) {real, imag} */,
  {32'h424685e8, 32'h42eeecde} /* (31, 10, 3) {real, imag} */,
  {32'hc327fb8b, 32'hc2ec3bea} /* (31, 10, 2) {real, imag} */,
  {32'h439c28bd, 32'hc23513fb} /* (31, 10, 1) {real, imag} */,
  {32'h416d1990, 32'h00000000} /* (31, 10, 0) {real, imag} */,
  {32'h4417dab0, 32'h3f896b58} /* (31, 9, 31) {real, imag} */,
  {32'hc394fea3, 32'h433faf52} /* (31, 9, 30) {real, imag} */,
  {32'h41e3d4bc, 32'hc1dc95f8} /* (31, 9, 29) {real, imag} */,
  {32'h42bd9902, 32'hc253f8bb} /* (31, 9, 28) {real, imag} */,
  {32'hc2086dd5, 32'hc0744b30} /* (31, 9, 27) {real, imag} */,
  {32'hc1df9fe4, 32'hc29ff680} /* (31, 9, 26) {real, imag} */,
  {32'hc0643630, 32'hc2f37c49} /* (31, 9, 25) {real, imag} */,
  {32'h4086b9c0, 32'hbf493f60} /* (31, 9, 24) {real, imag} */,
  {32'hc19f64b6, 32'h4223ac3c} /* (31, 9, 23) {real, imag} */,
  {32'hc02e6310, 32'h4149daea} /* (31, 9, 22) {real, imag} */,
  {32'hc2c1af58, 32'h40cc7540} /* (31, 9, 21) {real, imag} */,
  {32'hc25a9bad, 32'h4242e674} /* (31, 9, 20) {real, imag} */,
  {32'hc15d5714, 32'hc25a0603} /* (31, 9, 19) {real, imag} */,
  {32'hc257b514, 32'hc1d05dd4} /* (31, 9, 18) {real, imag} */,
  {32'hc1eb9c90, 32'h425479e3} /* (31, 9, 17) {real, imag} */,
  {32'h426d1ffb, 32'h00000000} /* (31, 9, 16) {real, imag} */,
  {32'hc1eb9c90, 32'hc25479e3} /* (31, 9, 15) {real, imag} */,
  {32'hc257b514, 32'h41d05dd4} /* (31, 9, 14) {real, imag} */,
  {32'hc15d5714, 32'h425a0603} /* (31, 9, 13) {real, imag} */,
  {32'hc25a9bad, 32'hc242e674} /* (31, 9, 12) {real, imag} */,
  {32'hc2c1af58, 32'hc0cc7540} /* (31, 9, 11) {real, imag} */,
  {32'hc02e6310, 32'hc149daea} /* (31, 9, 10) {real, imag} */,
  {32'hc19f64b6, 32'hc223ac3c} /* (31, 9, 9) {real, imag} */,
  {32'h4086b9c0, 32'h3f493f60} /* (31, 9, 8) {real, imag} */,
  {32'hc0643630, 32'h42f37c49} /* (31, 9, 7) {real, imag} */,
  {32'hc1df9fe4, 32'h429ff680} /* (31, 9, 6) {real, imag} */,
  {32'hc2086dd5, 32'h40744b30} /* (31, 9, 5) {real, imag} */,
  {32'h42bd9902, 32'h4253f8bb} /* (31, 9, 4) {real, imag} */,
  {32'h41e3d4bc, 32'h41dc95f8} /* (31, 9, 3) {real, imag} */,
  {32'hc394fea3, 32'hc33faf52} /* (31, 9, 2) {real, imag} */,
  {32'h4417dab0, 32'hbf896b58} /* (31, 9, 1) {real, imag} */,
  {32'h4383d4e4, 32'h00000000} /* (31, 9, 0) {real, imag} */,
  {32'h442d3502, 32'hc2855a40} /* (31, 8, 31) {real, imag} */,
  {32'hc3884ace, 32'h4306031d} /* (31, 8, 30) {real, imag} */,
  {32'hc2d83c42, 32'h41ed1920} /* (31, 8, 29) {real, imag} */,
  {32'h431f8efc, 32'hbd9a3800} /* (31, 8, 28) {real, imag} */,
  {32'hc11246e4, 32'h427d75ae} /* (31, 8, 27) {real, imag} */,
  {32'hc1bd5630, 32'hc22ff72a} /* (31, 8, 26) {real, imag} */,
  {32'h419e8002, 32'hbf757240} /* (31, 8, 25) {real, imag} */,
  {32'hc1e99202, 32'h4039f548} /* (31, 8, 24) {real, imag} */,
  {32'h41a63d22, 32'hc09850c0} /* (31, 8, 23) {real, imag} */,
  {32'h413c9e05, 32'hc0b43ac0} /* (31, 8, 22) {real, imag} */,
  {32'hc119c995, 32'h42b1731f} /* (31, 8, 21) {real, imag} */,
  {32'h41e2b162, 32'h4213b075} /* (31, 8, 20) {real, imag} */,
  {32'hc290598d, 32'hc23308ea} /* (31, 8, 19) {real, imag} */,
  {32'h41e06cc5, 32'hc18a73d9} /* (31, 8, 18) {real, imag} */,
  {32'h418f1238, 32'h4216d8c5} /* (31, 8, 17) {real, imag} */,
  {32'hc0801648, 32'h00000000} /* (31, 8, 16) {real, imag} */,
  {32'h418f1238, 32'hc216d8c5} /* (31, 8, 15) {real, imag} */,
  {32'h41e06cc5, 32'h418a73d9} /* (31, 8, 14) {real, imag} */,
  {32'hc290598d, 32'h423308ea} /* (31, 8, 13) {real, imag} */,
  {32'h41e2b162, 32'hc213b075} /* (31, 8, 12) {real, imag} */,
  {32'hc119c995, 32'hc2b1731f} /* (31, 8, 11) {real, imag} */,
  {32'h413c9e05, 32'h40b43ac0} /* (31, 8, 10) {real, imag} */,
  {32'h41a63d22, 32'h409850c0} /* (31, 8, 9) {real, imag} */,
  {32'hc1e99202, 32'hc039f548} /* (31, 8, 8) {real, imag} */,
  {32'h419e8002, 32'h3f757240} /* (31, 8, 7) {real, imag} */,
  {32'hc1bd5630, 32'h422ff72a} /* (31, 8, 6) {real, imag} */,
  {32'hc11246e4, 32'hc27d75ae} /* (31, 8, 5) {real, imag} */,
  {32'h431f8efc, 32'h3d9a3800} /* (31, 8, 4) {real, imag} */,
  {32'hc2d83c42, 32'hc1ed1920} /* (31, 8, 3) {real, imag} */,
  {32'hc3884ace, 32'hc306031d} /* (31, 8, 2) {real, imag} */,
  {32'h442d3502, 32'h42855a40} /* (31, 8, 1) {real, imag} */,
  {32'h436daba5, 32'h00000000} /* (31, 8, 0) {real, imag} */,
  {32'h44314943, 32'h41f8cc5a} /* (31, 7, 31) {real, imag} */,
  {32'hc32f94ab, 32'h434f9568} /* (31, 7, 30) {real, imag} */,
  {32'hc2b5fde2, 32'hc2cf2a6b} /* (31, 7, 29) {real, imag} */,
  {32'h4317e195, 32'hc21d9934} /* (31, 7, 28) {real, imag} */,
  {32'hc2701eb7, 32'hc1dfb0ea} /* (31, 7, 27) {real, imag} */,
  {32'hc2aa79bd, 32'h424a3a8a} /* (31, 7, 26) {real, imag} */,
  {32'h425770ba, 32'hc28e3a29} /* (31, 7, 25) {real, imag} */,
  {32'hc29b8c49, 32'hc1d0377a} /* (31, 7, 24) {real, imag} */,
  {32'hc19d2e8b, 32'hc227216a} /* (31, 7, 23) {real, imag} */,
  {32'h429686c6, 32'hc123364e} /* (31, 7, 22) {real, imag} */,
  {32'hc2d9e840, 32'h424f5f18} /* (31, 7, 21) {real, imag} */,
  {32'hc0eea6b8, 32'hc2477e28} /* (31, 7, 20) {real, imag} */,
  {32'h421658ec, 32'hc23d141c} /* (31, 7, 19) {real, imag} */,
  {32'h41e34c65, 32'h426ccdf4} /* (31, 7, 18) {real, imag} */,
  {32'hc0cb7b7c, 32'hc1b1c0ee} /* (31, 7, 17) {real, imag} */,
  {32'hc230ea48, 32'h00000000} /* (31, 7, 16) {real, imag} */,
  {32'hc0cb7b7c, 32'h41b1c0ee} /* (31, 7, 15) {real, imag} */,
  {32'h41e34c65, 32'hc26ccdf4} /* (31, 7, 14) {real, imag} */,
  {32'h421658ec, 32'h423d141c} /* (31, 7, 13) {real, imag} */,
  {32'hc0eea6b8, 32'h42477e28} /* (31, 7, 12) {real, imag} */,
  {32'hc2d9e840, 32'hc24f5f18} /* (31, 7, 11) {real, imag} */,
  {32'h429686c6, 32'h4123364e} /* (31, 7, 10) {real, imag} */,
  {32'hc19d2e8b, 32'h4227216a} /* (31, 7, 9) {real, imag} */,
  {32'hc29b8c49, 32'h41d0377a} /* (31, 7, 8) {real, imag} */,
  {32'h425770ba, 32'h428e3a29} /* (31, 7, 7) {real, imag} */,
  {32'hc2aa79bd, 32'hc24a3a8a} /* (31, 7, 6) {real, imag} */,
  {32'hc2701eb7, 32'h41dfb0ea} /* (31, 7, 5) {real, imag} */,
  {32'h4317e195, 32'h421d9934} /* (31, 7, 4) {real, imag} */,
  {32'hc2b5fde2, 32'h42cf2a6b} /* (31, 7, 3) {real, imag} */,
  {32'hc32f94ab, 32'hc34f9568} /* (31, 7, 2) {real, imag} */,
  {32'h44314943, 32'hc1f8cc5a} /* (31, 7, 1) {real, imag} */,
  {32'h4366fc68, 32'h00000000} /* (31, 7, 0) {real, imag} */,
  {32'h442e86e3, 32'h40e283c0} /* (31, 6, 31) {real, imag} */,
  {32'hc35185b1, 32'h439efc87} /* (31, 6, 30) {real, imag} */,
  {32'hc1a72718, 32'hc117c1e9} /* (31, 6, 29) {real, imag} */,
  {32'h429a43f9, 32'hc31d38e0} /* (31, 6, 28) {real, imag} */,
  {32'hbf10f6a0, 32'h4249fbf2} /* (31, 6, 27) {real, imag} */,
  {32'h3f253370, 32'h420156ab} /* (31, 6, 26) {real, imag} */,
  {32'hc18761f7, 32'h422f7a3d} /* (31, 6, 25) {real, imag} */,
  {32'hc19aaec6, 32'hc271de9b} /* (31, 6, 24) {real, imag} */,
  {32'h41c3aa06, 32'h41f06ccd} /* (31, 6, 23) {real, imag} */,
  {32'h42534466, 32'hc2ca02e2} /* (31, 6, 22) {real, imag} */,
  {32'hc2981455, 32'h42a2ab4d} /* (31, 6, 21) {real, imag} */,
  {32'hc1cb9d2c, 32'h40a1796c} /* (31, 6, 20) {real, imag} */,
  {32'hc24af628, 32'hc21758e3} /* (31, 6, 19) {real, imag} */,
  {32'hc252300c, 32'h42333400} /* (31, 6, 18) {real, imag} */,
  {32'hc2805340, 32'h404395ec} /* (31, 6, 17) {real, imag} */,
  {32'hc04877d4, 32'h00000000} /* (31, 6, 16) {real, imag} */,
  {32'hc2805340, 32'hc04395ec} /* (31, 6, 15) {real, imag} */,
  {32'hc252300c, 32'hc2333400} /* (31, 6, 14) {real, imag} */,
  {32'hc24af628, 32'h421758e3} /* (31, 6, 13) {real, imag} */,
  {32'hc1cb9d2c, 32'hc0a1796c} /* (31, 6, 12) {real, imag} */,
  {32'hc2981455, 32'hc2a2ab4d} /* (31, 6, 11) {real, imag} */,
  {32'h42534466, 32'h42ca02e2} /* (31, 6, 10) {real, imag} */,
  {32'h41c3aa06, 32'hc1f06ccd} /* (31, 6, 9) {real, imag} */,
  {32'hc19aaec6, 32'h4271de9b} /* (31, 6, 8) {real, imag} */,
  {32'hc18761f7, 32'hc22f7a3d} /* (31, 6, 7) {real, imag} */,
  {32'h3f253370, 32'hc20156ab} /* (31, 6, 6) {real, imag} */,
  {32'hbf10f6a0, 32'hc249fbf2} /* (31, 6, 5) {real, imag} */,
  {32'h429a43f9, 32'h431d38e0} /* (31, 6, 4) {real, imag} */,
  {32'hc1a72718, 32'h4117c1e9} /* (31, 6, 3) {real, imag} */,
  {32'hc35185b1, 32'hc39efc87} /* (31, 6, 2) {real, imag} */,
  {32'h442e86e3, 32'hc0e283c0} /* (31, 6, 1) {real, imag} */,
  {32'h43547bab, 32'h00000000} /* (31, 6, 0) {real, imag} */,
  {32'h44033409, 32'hc3940fde} /* (31, 5, 31) {real, imag} */,
  {32'hc28da6e8, 32'h43a0d2ac} /* (31, 5, 30) {real, imag} */,
  {32'hc21e39dc, 32'hc1704bfa} /* (31, 5, 29) {real, imag} */,
  {32'hc2a7b1d8, 32'hc2c2cdea} /* (31, 5, 28) {real, imag} */,
  {32'hc2580b96, 32'h41ecc8c2} /* (31, 5, 27) {real, imag} */,
  {32'hc1843058, 32'h425d9540} /* (31, 5, 26) {real, imag} */,
  {32'hc0693a98, 32'h420438ec} /* (31, 5, 25) {real, imag} */,
  {32'h41d51b0b, 32'hc2544fa6} /* (31, 5, 24) {real, imag} */,
  {32'h424f54b4, 32'h41cded5b} /* (31, 5, 23) {real, imag} */,
  {32'h4203cb56, 32'hc23e0972} /* (31, 5, 22) {real, imag} */,
  {32'h40bbb8c4, 32'h42071d18} /* (31, 5, 21) {real, imag} */,
  {32'hc2c8a0b0, 32'hc2367158} /* (31, 5, 20) {real, imag} */,
  {32'hc311f55c, 32'hc108ee46} /* (31, 5, 19) {real, imag} */,
  {32'hc26f1f65, 32'h4203678c} /* (31, 5, 18) {real, imag} */,
  {32'hc1575e90, 32'hc053ddc8} /* (31, 5, 17) {real, imag} */,
  {32'h3ec81140, 32'h00000000} /* (31, 5, 16) {real, imag} */,
  {32'hc1575e90, 32'h4053ddc8} /* (31, 5, 15) {real, imag} */,
  {32'hc26f1f65, 32'hc203678c} /* (31, 5, 14) {real, imag} */,
  {32'hc311f55c, 32'h4108ee46} /* (31, 5, 13) {real, imag} */,
  {32'hc2c8a0b0, 32'h42367158} /* (31, 5, 12) {real, imag} */,
  {32'h40bbb8c4, 32'hc2071d18} /* (31, 5, 11) {real, imag} */,
  {32'h4203cb56, 32'h423e0972} /* (31, 5, 10) {real, imag} */,
  {32'h424f54b4, 32'hc1cded5b} /* (31, 5, 9) {real, imag} */,
  {32'h41d51b0b, 32'h42544fa6} /* (31, 5, 8) {real, imag} */,
  {32'hc0693a98, 32'hc20438ec} /* (31, 5, 7) {real, imag} */,
  {32'hc1843058, 32'hc25d9540} /* (31, 5, 6) {real, imag} */,
  {32'hc2580b96, 32'hc1ecc8c2} /* (31, 5, 5) {real, imag} */,
  {32'hc2a7b1d8, 32'h42c2cdea} /* (31, 5, 4) {real, imag} */,
  {32'hc21e39dc, 32'h41704bfa} /* (31, 5, 3) {real, imag} */,
  {32'hc28da6e8, 32'hc3a0d2ac} /* (31, 5, 2) {real, imag} */,
  {32'h44033409, 32'h43940fde} /* (31, 5, 1) {real, imag} */,
  {32'h4333b76b, 32'h00000000} /* (31, 5, 0) {real, imag} */,
  {32'h43b779fe, 32'hc3bad384} /* (31, 4, 31) {real, imag} */,
  {32'h42853443, 32'h43b082e0} /* (31, 4, 30) {real, imag} */,
  {32'hc28091c8, 32'h415d027f} /* (31, 4, 29) {real, imag} */,
  {32'hc2143cb6, 32'h424f4477} /* (31, 4, 28) {real, imag} */,
  {32'h423ee722, 32'h42ab729c} /* (31, 4, 27) {real, imag} */,
  {32'h410206fc, 32'h4204cfab} /* (31, 4, 26) {real, imag} */,
  {32'h428ccf44, 32'hc2b12a30} /* (31, 4, 25) {real, imag} */,
  {32'h42812788, 32'h426e7827} /* (31, 4, 24) {real, imag} */,
  {32'hc22a4363, 32'h41a34481} /* (31, 4, 23) {real, imag} */,
  {32'hc134a8b6, 32'hc118d6f5} /* (31, 4, 22) {real, imag} */,
  {32'hc1fd9a5a, 32'hc1f3da20} /* (31, 4, 21) {real, imag} */,
  {32'hc1e60da6, 32'hc023e6b0} /* (31, 4, 20) {real, imag} */,
  {32'h41ca41b0, 32'hc2236add} /* (31, 4, 19) {real, imag} */,
  {32'hc01d0b28, 32'h42660c27} /* (31, 4, 18) {real, imag} */,
  {32'h40e1ced0, 32'h4193c1ec} /* (31, 4, 17) {real, imag} */,
  {32'h41ea2393, 32'h00000000} /* (31, 4, 16) {real, imag} */,
  {32'h40e1ced0, 32'hc193c1ec} /* (31, 4, 15) {real, imag} */,
  {32'hc01d0b28, 32'hc2660c27} /* (31, 4, 14) {real, imag} */,
  {32'h41ca41b0, 32'h42236add} /* (31, 4, 13) {real, imag} */,
  {32'hc1e60da6, 32'h4023e6b0} /* (31, 4, 12) {real, imag} */,
  {32'hc1fd9a5a, 32'h41f3da20} /* (31, 4, 11) {real, imag} */,
  {32'hc134a8b6, 32'h4118d6f5} /* (31, 4, 10) {real, imag} */,
  {32'hc22a4363, 32'hc1a34481} /* (31, 4, 9) {real, imag} */,
  {32'h42812788, 32'hc26e7827} /* (31, 4, 8) {real, imag} */,
  {32'h428ccf44, 32'h42b12a30} /* (31, 4, 7) {real, imag} */,
  {32'h410206fc, 32'hc204cfab} /* (31, 4, 6) {real, imag} */,
  {32'h423ee722, 32'hc2ab729c} /* (31, 4, 5) {real, imag} */,
  {32'hc2143cb6, 32'hc24f4477} /* (31, 4, 4) {real, imag} */,
  {32'hc28091c8, 32'hc15d027f} /* (31, 4, 3) {real, imag} */,
  {32'h42853443, 32'hc3b082e0} /* (31, 4, 2) {real, imag} */,
  {32'h43b779fe, 32'h43bad384} /* (31, 4, 1) {real, imag} */,
  {32'h417f47a0, 32'h00000000} /* (31, 4, 0) {real, imag} */,
  {32'h43b86f93, 32'hc410bf40} /* (31, 3, 31) {real, imag} */,
  {32'h4258eec0, 32'h43a6e63d} /* (31, 3, 30) {real, imag} */,
  {32'hc12d9784, 32'h419043ed} /* (31, 3, 29) {real, imag} */,
  {32'h41a6af94, 32'h428d7cb2} /* (31, 3, 28) {real, imag} */,
  {32'hc1587db8, 32'h422bd870} /* (31, 3, 27) {real, imag} */,
  {32'hc2832888, 32'h42467a26} /* (31, 3, 26) {real, imag} */,
  {32'hc228b3f7, 32'hc2111e32} /* (31, 3, 25) {real, imag} */,
  {32'h42440acc, 32'hc171269c} /* (31, 3, 24) {real, imag} */,
  {32'hc22c224a, 32'h4277678c} /* (31, 3, 23) {real, imag} */,
  {32'hc1a4ebc0, 32'hc17fdaa2} /* (31, 3, 22) {real, imag} */,
  {32'h409c6678, 32'h4188fc1f} /* (31, 3, 21) {real, imag} */,
  {32'hc273a3f7, 32'h429a8422} /* (31, 3, 20) {real, imag} */,
  {32'hc28b69fd, 32'hc0fc98b0} /* (31, 3, 19) {real, imag} */,
  {32'hc0b0ce3c, 32'hc10e9cba} /* (31, 3, 18) {real, imag} */,
  {32'h4204c3ae, 32'h41fa3e64} /* (31, 3, 17) {real, imag} */,
  {32'hc1d9016e, 32'h00000000} /* (31, 3, 16) {real, imag} */,
  {32'h4204c3ae, 32'hc1fa3e64} /* (31, 3, 15) {real, imag} */,
  {32'hc0b0ce3c, 32'h410e9cba} /* (31, 3, 14) {real, imag} */,
  {32'hc28b69fd, 32'h40fc98b0} /* (31, 3, 13) {real, imag} */,
  {32'hc273a3f7, 32'hc29a8422} /* (31, 3, 12) {real, imag} */,
  {32'h409c6678, 32'hc188fc1f} /* (31, 3, 11) {real, imag} */,
  {32'hc1a4ebc0, 32'h417fdaa2} /* (31, 3, 10) {real, imag} */,
  {32'hc22c224a, 32'hc277678c} /* (31, 3, 9) {real, imag} */,
  {32'h42440acc, 32'h4171269c} /* (31, 3, 8) {real, imag} */,
  {32'hc228b3f7, 32'h42111e32} /* (31, 3, 7) {real, imag} */,
  {32'hc2832888, 32'hc2467a26} /* (31, 3, 6) {real, imag} */,
  {32'hc1587db8, 32'hc22bd870} /* (31, 3, 5) {real, imag} */,
  {32'h41a6af94, 32'hc28d7cb2} /* (31, 3, 4) {real, imag} */,
  {32'hc12d9784, 32'hc19043ed} /* (31, 3, 3) {real, imag} */,
  {32'h4258eec0, 32'hc3a6e63d} /* (31, 3, 2) {real, imag} */,
  {32'h43b86f93, 32'h4410bf40} /* (31, 3, 1) {real, imag} */,
  {32'h41d2c748, 32'h00000000} /* (31, 3, 0) {real, imag} */,
  {32'h43976384, 32'hc40ceb74} /* (31, 2, 31) {real, imag} */,
  {32'h425aa314, 32'h43644774} /* (31, 2, 30) {real, imag} */,
  {32'h423a3c74, 32'h40b0d650} /* (31, 2, 29) {real, imag} */,
  {32'hc2a5a013, 32'h42ce1b3c} /* (31, 2, 28) {real, imag} */,
  {32'hc274df5d, 32'h42303bba} /* (31, 2, 27) {real, imag} */,
  {32'hc25aff7a, 32'hc283f549} /* (31, 2, 26) {real, imag} */,
  {32'hc1939c06, 32'hc29939d2} /* (31, 2, 25) {real, imag} */,
  {32'h3eda6200, 32'hc13f9d3d} /* (31, 2, 24) {real, imag} */,
  {32'hc20279fd, 32'hbf7d1140} /* (31, 2, 23) {real, imag} */,
  {32'h4147c3f0, 32'h429b7d8b} /* (31, 2, 22) {real, imag} */,
  {32'h4144f1e2, 32'hc1c9a0b2} /* (31, 2, 21) {real, imag} */,
  {32'h42a646fe, 32'h418c48ea} /* (31, 2, 20) {real, imag} */,
  {32'h417a2702, 32'hc12262ac} /* (31, 2, 19) {real, imag} */,
  {32'h413c0e34, 32'h40286990} /* (31, 2, 18) {real, imag} */,
  {32'hc25c94fa, 32'hc1629b26} /* (31, 2, 17) {real, imag} */,
  {32'h41969ebe, 32'h00000000} /* (31, 2, 16) {real, imag} */,
  {32'hc25c94fa, 32'h41629b26} /* (31, 2, 15) {real, imag} */,
  {32'h413c0e34, 32'hc0286990} /* (31, 2, 14) {real, imag} */,
  {32'h417a2702, 32'h412262ac} /* (31, 2, 13) {real, imag} */,
  {32'h42a646fe, 32'hc18c48ea} /* (31, 2, 12) {real, imag} */,
  {32'h4144f1e2, 32'h41c9a0b2} /* (31, 2, 11) {real, imag} */,
  {32'h4147c3f0, 32'hc29b7d8b} /* (31, 2, 10) {real, imag} */,
  {32'hc20279fd, 32'h3f7d1140} /* (31, 2, 9) {real, imag} */,
  {32'h3eda6200, 32'h413f9d3d} /* (31, 2, 8) {real, imag} */,
  {32'hc1939c06, 32'h429939d2} /* (31, 2, 7) {real, imag} */,
  {32'hc25aff7a, 32'h4283f549} /* (31, 2, 6) {real, imag} */,
  {32'hc274df5d, 32'hc2303bba} /* (31, 2, 5) {real, imag} */,
  {32'hc2a5a013, 32'hc2ce1b3c} /* (31, 2, 4) {real, imag} */,
  {32'h423a3c74, 32'hc0b0d650} /* (31, 2, 3) {real, imag} */,
  {32'h425aa314, 32'hc3644774} /* (31, 2, 2) {real, imag} */,
  {32'h43976384, 32'h440ceb74} /* (31, 2, 1) {real, imag} */,
  {32'hc28c2bbc, 32'h00000000} /* (31, 2, 0) {real, imag} */,
  {32'h4343ede6, 32'hc3fdeb9c} /* (31, 1, 31) {real, imag} */,
  {32'hc1bd7c78, 32'h434083a6} /* (31, 1, 30) {real, imag} */,
  {32'hc118b13e, 32'h42d2f07a} /* (31, 1, 29) {real, imag} */,
  {32'hc29cd22a, 32'h422c0aff} /* (31, 1, 28) {real, imag} */,
  {32'h413d355c, 32'hc137e025} /* (31, 1, 27) {real, imag} */,
  {32'hc28049b3, 32'hbf09cde0} /* (31, 1, 26) {real, imag} */,
  {32'hbfde7520, 32'hc29488d0} /* (31, 1, 25) {real, imag} */,
  {32'h428c3575, 32'h40de2b80} /* (31, 1, 24) {real, imag} */,
  {32'hc28ae470, 32'hc2163c86} /* (31, 1, 23) {real, imag} */,
  {32'hc29032a7, 32'h409dc2f6} /* (31, 1, 22) {real, imag} */,
  {32'hc239d714, 32'h419caa4e} /* (31, 1, 21) {real, imag} */,
  {32'h4241d148, 32'hc1363e36} /* (31, 1, 20) {real, imag} */,
  {32'h4227035e, 32'h40035abc} /* (31, 1, 19) {real, imag} */,
  {32'h41244143, 32'hc10dc19d} /* (31, 1, 18) {real, imag} */,
  {32'h4175773e, 32'h4293f625} /* (31, 1, 17) {real, imag} */,
  {32'hc1ae9903, 32'h00000000} /* (31, 1, 16) {real, imag} */,
  {32'h4175773e, 32'hc293f625} /* (31, 1, 15) {real, imag} */,
  {32'h41244143, 32'h410dc19d} /* (31, 1, 14) {real, imag} */,
  {32'h4227035e, 32'hc0035abc} /* (31, 1, 13) {real, imag} */,
  {32'h4241d148, 32'h41363e36} /* (31, 1, 12) {real, imag} */,
  {32'hc239d714, 32'hc19caa4e} /* (31, 1, 11) {real, imag} */,
  {32'hc29032a7, 32'hc09dc2f6} /* (31, 1, 10) {real, imag} */,
  {32'hc28ae470, 32'h42163c86} /* (31, 1, 9) {real, imag} */,
  {32'h428c3575, 32'hc0de2b80} /* (31, 1, 8) {real, imag} */,
  {32'hbfde7520, 32'h429488d0} /* (31, 1, 7) {real, imag} */,
  {32'hc28049b3, 32'h3f09cde0} /* (31, 1, 6) {real, imag} */,
  {32'h413d355c, 32'h4137e025} /* (31, 1, 5) {real, imag} */,
  {32'hc29cd22a, 32'hc22c0aff} /* (31, 1, 4) {real, imag} */,
  {32'hc118b13e, 32'hc2d2f07a} /* (31, 1, 3) {real, imag} */,
  {32'hc1bd7c78, 32'hc34083a6} /* (31, 1, 2) {real, imag} */,
  {32'h4343ede6, 32'h43fdeb9c} /* (31, 1, 1) {real, imag} */,
  {32'h41e35728, 32'h00000000} /* (31, 1, 0) {real, imag} */,
  {32'h433dd736, 32'hc3b2f0e7} /* (31, 0, 31) {real, imag} */,
  {32'hc30d5d50, 32'h43740a7f} /* (31, 0, 30) {real, imag} */,
  {32'h41d25d5e, 32'h41656708} /* (31, 0, 29) {real, imag} */,
  {32'hc0745fc0, 32'h41e884d8} /* (31, 0, 28) {real, imag} */,
  {32'h407caa70, 32'hc24384ae} /* (31, 0, 27) {real, imag} */,
  {32'h41110580, 32'h41328b12} /* (31, 0, 26) {real, imag} */,
  {32'hc1c226a0, 32'hc1e6f212} /* (31, 0, 25) {real, imag} */,
  {32'h41cef778, 32'hbec45180} /* (31, 0, 24) {real, imag} */,
  {32'hc1abcd3d, 32'h41fc0f38} /* (31, 0, 23) {real, imag} */,
  {32'h41c1d12a, 32'hc152b8e6} /* (31, 0, 22) {real, imag} */,
  {32'hc0b17a90, 32'hc198b946} /* (31, 0, 21) {real, imag} */,
  {32'hc1c1e548, 32'h4211d5c3} /* (31, 0, 20) {real, imag} */,
  {32'hc234dfe5, 32'hc1df0776} /* (31, 0, 19) {real, imag} */,
  {32'h41c255f6, 32'hc1e8c622} /* (31, 0, 18) {real, imag} */,
  {32'h41423924, 32'h4022b2f4} /* (31, 0, 17) {real, imag} */,
  {32'hc1e6bf08, 32'h00000000} /* (31, 0, 16) {real, imag} */,
  {32'h41423924, 32'hc022b2f4} /* (31, 0, 15) {real, imag} */,
  {32'h41c255f6, 32'h41e8c622} /* (31, 0, 14) {real, imag} */,
  {32'hc234dfe5, 32'h41df0776} /* (31, 0, 13) {real, imag} */,
  {32'hc1c1e548, 32'hc211d5c3} /* (31, 0, 12) {real, imag} */,
  {32'hc0b17a90, 32'h4198b946} /* (31, 0, 11) {real, imag} */,
  {32'h41c1d12a, 32'h4152b8e6} /* (31, 0, 10) {real, imag} */,
  {32'hc1abcd3d, 32'hc1fc0f38} /* (31, 0, 9) {real, imag} */,
  {32'h41cef778, 32'h3ec45180} /* (31, 0, 8) {real, imag} */,
  {32'hc1c226a0, 32'h41e6f212} /* (31, 0, 7) {real, imag} */,
  {32'h41110580, 32'hc1328b12} /* (31, 0, 6) {real, imag} */,
  {32'h407caa70, 32'h424384ae} /* (31, 0, 5) {real, imag} */,
  {32'hc0745fc0, 32'hc1e884d8} /* (31, 0, 4) {real, imag} */,
  {32'h41d25d5e, 32'hc1656708} /* (31, 0, 3) {real, imag} */,
  {32'hc30d5d50, 32'hc3740a7f} /* (31, 0, 2) {real, imag} */,
  {32'h433dd736, 32'h43b2f0e7} /* (31, 0, 1) {real, imag} */,
  {32'h420bf0bc, 32'h00000000} /* (31, 0, 0) {real, imag} */,
  {32'h445624b8, 32'hc40cac78} /* (30, 31, 31) {real, imag} */,
  {32'hc3c0a9ae, 32'h43d10372} /* (30, 31, 30) {real, imag} */,
  {32'hc1f5ab1c, 32'hc1fa3e90} /* (30, 31, 29) {real, imag} */,
  {32'h42d4afe9, 32'h427de6f2} /* (30, 31, 28) {real, imag} */,
  {32'hc2994eff, 32'h41daa400} /* (30, 31, 27) {real, imag} */,
  {32'hc24dab27, 32'hc22f5398} /* (30, 31, 26) {real, imag} */,
  {32'hc16f07bc, 32'h4220410e} /* (30, 31, 25) {real, imag} */,
  {32'hc0f9e95c, 32'h42cf2593} /* (30, 31, 24) {real, imag} */,
  {32'h429f4969, 32'h4126b794} /* (30, 31, 23) {real, imag} */,
  {32'hc23fed74, 32'hc290c04b} /* (30, 31, 22) {real, imag} */,
  {32'hc0d36408, 32'h410e1ddc} /* (30, 31, 21) {real, imag} */,
  {32'hc0c19da9, 32'h41101b4e} /* (30, 31, 20) {real, imag} */,
  {32'h4232acb4, 32'h40c75390} /* (30, 31, 19) {real, imag} */,
  {32'h40dd3f42, 32'hc1930e86} /* (30, 31, 18) {real, imag} */,
  {32'hc0c4bd6c, 32'hc2957000} /* (30, 31, 17) {real, imag} */,
  {32'hc22df4c2, 32'h00000000} /* (30, 31, 16) {real, imag} */,
  {32'hc0c4bd6c, 32'h42957000} /* (30, 31, 15) {real, imag} */,
  {32'h40dd3f42, 32'h41930e86} /* (30, 31, 14) {real, imag} */,
  {32'h4232acb4, 32'hc0c75390} /* (30, 31, 13) {real, imag} */,
  {32'hc0c19da9, 32'hc1101b4e} /* (30, 31, 12) {real, imag} */,
  {32'hc0d36408, 32'hc10e1ddc} /* (30, 31, 11) {real, imag} */,
  {32'hc23fed74, 32'h4290c04b} /* (30, 31, 10) {real, imag} */,
  {32'h429f4969, 32'hc126b794} /* (30, 31, 9) {real, imag} */,
  {32'hc0f9e95c, 32'hc2cf2593} /* (30, 31, 8) {real, imag} */,
  {32'hc16f07bc, 32'hc220410e} /* (30, 31, 7) {real, imag} */,
  {32'hc24dab27, 32'h422f5398} /* (30, 31, 6) {real, imag} */,
  {32'hc2994eff, 32'hc1daa400} /* (30, 31, 5) {real, imag} */,
  {32'h42d4afe9, 32'hc27de6f2} /* (30, 31, 4) {real, imag} */,
  {32'hc1f5ab1c, 32'h41fa3e90} /* (30, 31, 3) {real, imag} */,
  {32'hc3c0a9ae, 32'hc3d10372} /* (30, 31, 2) {real, imag} */,
  {32'h445624b8, 32'h440cac78} /* (30, 31, 1) {real, imag} */,
  {32'h43d265ae, 32'h00000000} /* (30, 31, 0) {real, imag} */,
  {32'h44a64438, 32'hc40eff1e} /* (30, 30, 31) {real, imag} */,
  {32'hc4314c4e, 32'h44060756} /* (30, 30, 30) {real, imag} */,
  {32'h41e543ea, 32'hc2663d78} /* (30, 30, 29) {real, imag} */,
  {32'h43695a64, 32'h42b09ae0} /* (30, 30, 28) {real, imag} */,
  {32'hc340ded8, 32'h41b12f50} /* (30, 30, 27) {real, imag} */,
  {32'h428fe00c, 32'hc31cced5} /* (30, 30, 26) {real, imag} */,
  {32'hc20bedfa, 32'h428aa031} /* (30, 30, 25) {real, imag} */,
  {32'h42222345, 32'h42b9f86c} /* (30, 30, 24) {real, imag} */,
  {32'h4282747a, 32'h429d3a4c} /* (30, 30, 23) {real, imag} */,
  {32'hc21319a8, 32'h42361605} /* (30, 30, 22) {real, imag} */,
  {32'h42001fc9, 32'h4251cc5a} /* (30, 30, 21) {real, imag} */,
  {32'h408dd968, 32'h4226b26e} /* (30, 30, 20) {real, imag} */,
  {32'hc2588896, 32'h411dfcb6} /* (30, 30, 19) {real, imag} */,
  {32'h414d23c8, 32'h4208e225} /* (30, 30, 18) {real, imag} */,
  {32'hc01186d8, 32'hc26ca192} /* (30, 30, 17) {real, imag} */,
  {32'hc12c6958, 32'h00000000} /* (30, 30, 16) {real, imag} */,
  {32'hc01186d8, 32'h426ca192} /* (30, 30, 15) {real, imag} */,
  {32'h414d23c8, 32'hc208e225} /* (30, 30, 14) {real, imag} */,
  {32'hc2588896, 32'hc11dfcb6} /* (30, 30, 13) {real, imag} */,
  {32'h408dd968, 32'hc226b26e} /* (30, 30, 12) {real, imag} */,
  {32'h42001fc9, 32'hc251cc5a} /* (30, 30, 11) {real, imag} */,
  {32'hc21319a8, 32'hc2361605} /* (30, 30, 10) {real, imag} */,
  {32'h4282747a, 32'hc29d3a4c} /* (30, 30, 9) {real, imag} */,
  {32'h42222345, 32'hc2b9f86c} /* (30, 30, 8) {real, imag} */,
  {32'hc20bedfa, 32'hc28aa031} /* (30, 30, 7) {real, imag} */,
  {32'h428fe00c, 32'h431cced5} /* (30, 30, 6) {real, imag} */,
  {32'hc340ded8, 32'hc1b12f50} /* (30, 30, 5) {real, imag} */,
  {32'h43695a64, 32'hc2b09ae0} /* (30, 30, 4) {real, imag} */,
  {32'h41e543ea, 32'h42663d78} /* (30, 30, 3) {real, imag} */,
  {32'hc4314c4e, 32'hc4060756} /* (30, 30, 2) {real, imag} */,
  {32'h44a64438, 32'h440eff1e} /* (30, 30, 1) {real, imag} */,
  {32'h4441eb6e, 32'h00000000} /* (30, 30, 0) {real, imag} */,
  {32'h44b27294, 32'hc3ab1f66} /* (30, 29, 31) {real, imag} */,
  {32'hc44a9b09, 32'h43ca0e2c} /* (30, 29, 30) {real, imag} */,
  {32'h41043560, 32'hc1f2ac4c} /* (30, 29, 29) {real, imag} */,
  {32'h431015e2, 32'hc1b29fc8} /* (30, 29, 28) {real, imag} */,
  {32'hc35d6993, 32'hc1fc72a6} /* (30, 29, 27) {real, imag} */,
  {32'hc301668f, 32'hc1c06f08} /* (30, 29, 26) {real, imag} */,
  {32'h42829348, 32'hc200b666} /* (30, 29, 25) {real, imag} */,
  {32'hc1d04004, 32'h42892f58} /* (30, 29, 24) {real, imag} */,
  {32'h41aa0c06, 32'h4226195c} /* (30, 29, 23) {real, imag} */,
  {32'hc1bad18d, 32'hc2ae23e9} /* (30, 29, 22) {real, imag} */,
  {32'h42756f21, 32'h4269e3c2} /* (30, 29, 21) {real, imag} */,
  {32'h425a035c, 32'h42648ca7} /* (30, 29, 20) {real, imag} */,
  {32'h428cc015, 32'h4076adb0} /* (30, 29, 19) {real, imag} */,
  {32'hc0fdee6c, 32'h421578da} /* (30, 29, 18) {real, imag} */,
  {32'h418fdc81, 32'h42698c0a} /* (30, 29, 17) {real, imag} */,
  {32'hc2a9610a, 32'h00000000} /* (30, 29, 16) {real, imag} */,
  {32'h418fdc81, 32'hc2698c0a} /* (30, 29, 15) {real, imag} */,
  {32'hc0fdee6c, 32'hc21578da} /* (30, 29, 14) {real, imag} */,
  {32'h428cc015, 32'hc076adb0} /* (30, 29, 13) {real, imag} */,
  {32'h425a035c, 32'hc2648ca7} /* (30, 29, 12) {real, imag} */,
  {32'h42756f21, 32'hc269e3c2} /* (30, 29, 11) {real, imag} */,
  {32'hc1bad18d, 32'h42ae23e9} /* (30, 29, 10) {real, imag} */,
  {32'h41aa0c06, 32'hc226195c} /* (30, 29, 9) {real, imag} */,
  {32'hc1d04004, 32'hc2892f58} /* (30, 29, 8) {real, imag} */,
  {32'h42829348, 32'h4200b666} /* (30, 29, 7) {real, imag} */,
  {32'hc301668f, 32'h41c06f08} /* (30, 29, 6) {real, imag} */,
  {32'hc35d6993, 32'h41fc72a6} /* (30, 29, 5) {real, imag} */,
  {32'h431015e2, 32'h41b29fc8} /* (30, 29, 4) {real, imag} */,
  {32'h41043560, 32'h41f2ac4c} /* (30, 29, 3) {real, imag} */,
  {32'hc44a9b09, 32'hc3ca0e2c} /* (30, 29, 2) {real, imag} */,
  {32'h44b27294, 32'h43ab1f66} /* (30, 29, 1) {real, imag} */,
  {32'h441dc60c, 32'h00000000} /* (30, 29, 0) {real, imag} */,
  {32'h44b89d90, 32'hc3363c34} /* (30, 28, 31) {real, imag} */,
  {32'hc44d50fb, 32'h42bc00ac} /* (30, 28, 30) {real, imag} */,
  {32'hc30bbb30, 32'hc2a19154} /* (30, 28, 29) {real, imag} */,
  {32'h43228b48, 32'hc204b56a} /* (30, 28, 28) {real, imag} */,
  {32'hc3314d84, 32'hc1f79cc8} /* (30, 28, 27) {real, imag} */,
  {32'hc271209a, 32'hc063e038} /* (30, 28, 26) {real, imag} */,
  {32'hc3002bce, 32'hc21162ba} /* (30, 28, 25) {real, imag} */,
  {32'hc2941b51, 32'h42c36309} /* (30, 28, 24) {real, imag} */,
  {32'hc0603cac, 32'h42e5bfa6} /* (30, 28, 23) {real, imag} */,
  {32'h424149d1, 32'hc1216a77} /* (30, 28, 22) {real, imag} */,
  {32'h42c5a306, 32'h42a23fb8} /* (30, 28, 21) {real, imag} */,
  {32'h4292e1a8, 32'hc1bca943} /* (30, 28, 20) {real, imag} */,
  {32'h420d89a4, 32'h4181b992} /* (30, 28, 19) {real, imag} */,
  {32'hc28651f7, 32'hc1430ebc} /* (30, 28, 18) {real, imag} */,
  {32'h3e8a7500, 32'hc28b06ac} /* (30, 28, 17) {real, imag} */,
  {32'h42674c33, 32'h00000000} /* (30, 28, 16) {real, imag} */,
  {32'h3e8a7500, 32'h428b06ac} /* (30, 28, 15) {real, imag} */,
  {32'hc28651f7, 32'h41430ebc} /* (30, 28, 14) {real, imag} */,
  {32'h420d89a4, 32'hc181b992} /* (30, 28, 13) {real, imag} */,
  {32'h4292e1a8, 32'h41bca943} /* (30, 28, 12) {real, imag} */,
  {32'h42c5a306, 32'hc2a23fb8} /* (30, 28, 11) {real, imag} */,
  {32'h424149d1, 32'h41216a77} /* (30, 28, 10) {real, imag} */,
  {32'hc0603cac, 32'hc2e5bfa6} /* (30, 28, 9) {real, imag} */,
  {32'hc2941b51, 32'hc2c36309} /* (30, 28, 8) {real, imag} */,
  {32'hc3002bce, 32'h421162ba} /* (30, 28, 7) {real, imag} */,
  {32'hc271209a, 32'h4063e038} /* (30, 28, 6) {real, imag} */,
  {32'hc3314d84, 32'h41f79cc8} /* (30, 28, 5) {real, imag} */,
  {32'h43228b48, 32'h4204b56a} /* (30, 28, 4) {real, imag} */,
  {32'hc30bbb30, 32'h42a19154} /* (30, 28, 3) {real, imag} */,
  {32'hc44d50fb, 32'hc2bc00ac} /* (30, 28, 2) {real, imag} */,
  {32'h44b89d90, 32'h43363c34} /* (30, 28, 1) {real, imag} */,
  {32'h44419a58, 32'h00000000} /* (30, 28, 0) {real, imag} */,
  {32'h44b39a36, 32'hc2e1cfb0} /* (30, 27, 31) {real, imag} */,
  {32'hc4746f7c, 32'h43439905} /* (30, 27, 30) {real, imag} */,
  {32'hc15faad4, 32'hc3408951} /* (30, 27, 29) {real, imag} */,
  {32'h431c5eb6, 32'h42bfdb68} /* (30, 27, 28) {real, imag} */,
  {32'hc2e7ba5e, 32'h42733baa} /* (30, 27, 27) {real, imag} */,
  {32'h42738a19, 32'hc308b7ea} /* (30, 27, 26) {real, imag} */,
  {32'hc2dde7a1, 32'hc302871d} /* (30, 27, 25) {real, imag} */,
  {32'hc21ad470, 32'h42488a38} /* (30, 27, 24) {real, imag} */,
  {32'hc282918e, 32'h42921f76} /* (30, 27, 23) {real, imag} */,
  {32'h42384c1e, 32'hc10a4534} /* (30, 27, 22) {real, imag} */,
  {32'h424941a0, 32'h427a384d} /* (30, 27, 21) {real, imag} */,
  {32'hc2df6850, 32'hc24f1772} /* (30, 27, 20) {real, imag} */,
  {32'hc200e04a, 32'hc3036b8c} /* (30, 27, 19) {real, imag} */,
  {32'hc0d3e6f5, 32'h429e8bd0} /* (30, 27, 18) {real, imag} */,
  {32'hc1f13533, 32'hc202d879} /* (30, 27, 17) {real, imag} */,
  {32'h41b7ac4e, 32'h00000000} /* (30, 27, 16) {real, imag} */,
  {32'hc1f13533, 32'h4202d879} /* (30, 27, 15) {real, imag} */,
  {32'hc0d3e6f5, 32'hc29e8bd0} /* (30, 27, 14) {real, imag} */,
  {32'hc200e04a, 32'h43036b8c} /* (30, 27, 13) {real, imag} */,
  {32'hc2df6850, 32'h424f1772} /* (30, 27, 12) {real, imag} */,
  {32'h424941a0, 32'hc27a384d} /* (30, 27, 11) {real, imag} */,
  {32'h42384c1e, 32'h410a4534} /* (30, 27, 10) {real, imag} */,
  {32'hc282918e, 32'hc2921f76} /* (30, 27, 9) {real, imag} */,
  {32'hc21ad470, 32'hc2488a38} /* (30, 27, 8) {real, imag} */,
  {32'hc2dde7a1, 32'h4302871d} /* (30, 27, 7) {real, imag} */,
  {32'h42738a19, 32'h4308b7ea} /* (30, 27, 6) {real, imag} */,
  {32'hc2e7ba5e, 32'hc2733baa} /* (30, 27, 5) {real, imag} */,
  {32'h431c5eb6, 32'hc2bfdb68} /* (30, 27, 4) {real, imag} */,
  {32'hc15faad4, 32'h43408951} /* (30, 27, 3) {real, imag} */,
  {32'hc4746f7c, 32'hc3439905} /* (30, 27, 2) {real, imag} */,
  {32'h44b39a36, 32'h42e1cfb0} /* (30, 27, 1) {real, imag} */,
  {32'h44761818, 32'h00000000} /* (30, 27, 0) {real, imag} */,
  {32'h44bae5d8, 32'hc29ac036} /* (30, 26, 31) {real, imag} */,
  {32'hc45ece16, 32'h43ab95be} /* (30, 26, 30) {real, imag} */,
  {32'hc2bce90a, 32'hc2e2032a} /* (30, 26, 29) {real, imag} */,
  {32'h432a57f5, 32'h424dae6f} /* (30, 26, 28) {real, imag} */,
  {32'hc2d5ac3a, 32'h427951de} /* (30, 26, 27) {real, imag} */,
  {32'hc2747ca9, 32'h422b8fce} /* (30, 26, 26) {real, imag} */,
  {32'hc29bbb6c, 32'hc2889d38} /* (30, 26, 25) {real, imag} */,
  {32'hc2a0ca5e, 32'h425b3ae5} /* (30, 26, 24) {real, imag} */,
  {32'hc0230f50, 32'hc2c3a7bd} /* (30, 26, 23) {real, imag} */,
  {32'h4128c010, 32'hc1f55170} /* (30, 26, 22) {real, imag} */,
  {32'h41a37152, 32'h424b48ba} /* (30, 26, 21) {real, imag} */,
  {32'h42b34b96, 32'h42483664} /* (30, 26, 20) {real, imag} */,
  {32'h4194fe73, 32'hbfd495b0} /* (30, 26, 19) {real, imag} */,
  {32'h41b2adaf, 32'hc05490b0} /* (30, 26, 18) {real, imag} */,
  {32'hc21b6602, 32'hc0eaac8c} /* (30, 26, 17) {real, imag} */,
  {32'hbe40dd00, 32'h00000000} /* (30, 26, 16) {real, imag} */,
  {32'hc21b6602, 32'h40eaac8c} /* (30, 26, 15) {real, imag} */,
  {32'h41b2adaf, 32'h405490b0} /* (30, 26, 14) {real, imag} */,
  {32'h4194fe73, 32'h3fd495b0} /* (30, 26, 13) {real, imag} */,
  {32'h42b34b96, 32'hc2483664} /* (30, 26, 12) {real, imag} */,
  {32'h41a37152, 32'hc24b48ba} /* (30, 26, 11) {real, imag} */,
  {32'h4128c010, 32'h41f55170} /* (30, 26, 10) {real, imag} */,
  {32'hc0230f50, 32'h42c3a7bd} /* (30, 26, 9) {real, imag} */,
  {32'hc2a0ca5e, 32'hc25b3ae5} /* (30, 26, 8) {real, imag} */,
  {32'hc29bbb6c, 32'h42889d38} /* (30, 26, 7) {real, imag} */,
  {32'hc2747ca9, 32'hc22b8fce} /* (30, 26, 6) {real, imag} */,
  {32'hc2d5ac3a, 32'hc27951de} /* (30, 26, 5) {real, imag} */,
  {32'h432a57f5, 32'hc24dae6f} /* (30, 26, 4) {real, imag} */,
  {32'hc2bce90a, 32'h42e2032a} /* (30, 26, 3) {real, imag} */,
  {32'hc45ece16, 32'hc3ab95be} /* (30, 26, 2) {real, imag} */,
  {32'h44bae5d8, 32'h429ac036} /* (30, 26, 1) {real, imag} */,
  {32'h4473b27c, 32'h00000000} /* (30, 26, 0) {real, imag} */,
  {32'h44c5e649, 32'hc2b0a720} /* (30, 25, 31) {real, imag} */,
  {32'hc48527fa, 32'h438c7e20} /* (30, 25, 30) {real, imag} */,
  {32'hc2d89c4c, 32'hc2dea51a} /* (30, 25, 29) {real, imag} */,
  {32'h428aa9e4, 32'h411aec16} /* (30, 25, 28) {real, imag} */,
  {32'hc315fb2d, 32'hc2277855} /* (30, 25, 27) {real, imag} */,
  {32'h4248d6ac, 32'hc2abed6a} /* (30, 25, 26) {real, imag} */,
  {32'hc23b676e, 32'hc2b7b7be} /* (30, 25, 25) {real, imag} */,
  {32'hc2b1a3e8, 32'h41ab049d} /* (30, 25, 24) {real, imag} */,
  {32'h3fb56398, 32'h4251a807} /* (30, 25, 23) {real, imag} */,
  {32'hc2a5914c, 32'hc0fda338} /* (30, 25, 22) {real, imag} */,
  {32'hc2861006, 32'h42f39d01} /* (30, 25, 21) {real, imag} */,
  {32'h428c88ac, 32'hc2a2145b} /* (30, 25, 20) {real, imag} */,
  {32'h426bc3b0, 32'h42714b68} /* (30, 25, 19) {real, imag} */,
  {32'h41d67c1a, 32'hc137adac} /* (30, 25, 18) {real, imag} */,
  {32'h41e89787, 32'hc1bcc8aa} /* (30, 25, 17) {real, imag} */,
  {32'hc1e9c721, 32'h00000000} /* (30, 25, 16) {real, imag} */,
  {32'h41e89787, 32'h41bcc8aa} /* (30, 25, 15) {real, imag} */,
  {32'h41d67c1a, 32'h4137adac} /* (30, 25, 14) {real, imag} */,
  {32'h426bc3b0, 32'hc2714b68} /* (30, 25, 13) {real, imag} */,
  {32'h428c88ac, 32'h42a2145b} /* (30, 25, 12) {real, imag} */,
  {32'hc2861006, 32'hc2f39d01} /* (30, 25, 11) {real, imag} */,
  {32'hc2a5914c, 32'h40fda338} /* (30, 25, 10) {real, imag} */,
  {32'h3fb56398, 32'hc251a807} /* (30, 25, 9) {real, imag} */,
  {32'hc2b1a3e8, 32'hc1ab049d} /* (30, 25, 8) {real, imag} */,
  {32'hc23b676e, 32'h42b7b7be} /* (30, 25, 7) {real, imag} */,
  {32'h4248d6ac, 32'h42abed6a} /* (30, 25, 6) {real, imag} */,
  {32'hc315fb2d, 32'h42277855} /* (30, 25, 5) {real, imag} */,
  {32'h428aa9e4, 32'hc11aec16} /* (30, 25, 4) {real, imag} */,
  {32'hc2d89c4c, 32'h42dea51a} /* (30, 25, 3) {real, imag} */,
  {32'hc48527fa, 32'hc38c7e20} /* (30, 25, 2) {real, imag} */,
  {32'h44c5e649, 32'h42b0a720} /* (30, 25, 1) {real, imag} */,
  {32'h44618a60, 32'h00000000} /* (30, 25, 0) {real, imag} */,
  {32'h44b710d6, 32'h42446ea4} /* (30, 24, 31) {real, imag} */,
  {32'hc457c692, 32'h43985608} /* (30, 24, 30) {real, imag} */,
  {32'h4122eaa0, 32'hc26725aa} /* (30, 24, 29) {real, imag} */,
  {32'h42993f12, 32'hc2d4d546} /* (30, 24, 28) {real, imag} */,
  {32'hc34c97a6, 32'hc0392ad0} /* (30, 24, 27) {real, imag} */,
  {32'hc29fc565, 32'h41664f5c} /* (30, 24, 26) {real, imag} */,
  {32'hc2b61439, 32'hc2ea34ec} /* (30, 24, 25) {real, imag} */,
  {32'hc30fdbb3, 32'h422f3fc9} /* (30, 24, 24) {real, imag} */,
  {32'h41a09de4, 32'h4301fa1e} /* (30, 24, 23) {real, imag} */,
  {32'h41882ab4, 32'hc3014db3} /* (30, 24, 22) {real, imag} */,
  {32'h420012ea, 32'hc1aa5da6} /* (30, 24, 21) {real, imag} */,
  {32'h41bf88c2, 32'hc2c3be31} /* (30, 24, 20) {real, imag} */,
  {32'hc1673f44, 32'hc21e1e57} /* (30, 24, 19) {real, imag} */,
  {32'hc1c47aac, 32'h42d80608} /* (30, 24, 18) {real, imag} */,
  {32'h41460b54, 32'h42005377} /* (30, 24, 17) {real, imag} */,
  {32'hc2013bb8, 32'h00000000} /* (30, 24, 16) {real, imag} */,
  {32'h41460b54, 32'hc2005377} /* (30, 24, 15) {real, imag} */,
  {32'hc1c47aac, 32'hc2d80608} /* (30, 24, 14) {real, imag} */,
  {32'hc1673f44, 32'h421e1e57} /* (30, 24, 13) {real, imag} */,
  {32'h41bf88c2, 32'h42c3be31} /* (30, 24, 12) {real, imag} */,
  {32'h420012ea, 32'h41aa5da6} /* (30, 24, 11) {real, imag} */,
  {32'h41882ab4, 32'h43014db3} /* (30, 24, 10) {real, imag} */,
  {32'h41a09de4, 32'hc301fa1e} /* (30, 24, 9) {real, imag} */,
  {32'hc30fdbb3, 32'hc22f3fc9} /* (30, 24, 8) {real, imag} */,
  {32'hc2b61439, 32'h42ea34ec} /* (30, 24, 7) {real, imag} */,
  {32'hc29fc565, 32'hc1664f5c} /* (30, 24, 6) {real, imag} */,
  {32'hc34c97a6, 32'h40392ad0} /* (30, 24, 5) {real, imag} */,
  {32'h42993f12, 32'h42d4d546} /* (30, 24, 4) {real, imag} */,
  {32'h4122eaa0, 32'h426725aa} /* (30, 24, 3) {real, imag} */,
  {32'hc457c692, 32'hc3985608} /* (30, 24, 2) {real, imag} */,
  {32'h44b710d6, 32'hc2446ea4} /* (30, 24, 1) {real, imag} */,
  {32'h447c3498, 32'h00000000} /* (30, 24, 0) {real, imag} */,
  {32'h449257fa, 32'h42866420} /* (30, 23, 31) {real, imag} */,
  {32'hc4258a3f, 32'h43a6be8b} /* (30, 23, 30) {real, imag} */,
  {32'h4318d446, 32'h422536c8} /* (30, 23, 29) {real, imag} */,
  {32'h42d78c41, 32'hc2e43a0a} /* (30, 23, 28) {real, imag} */,
  {32'hc31a834e, 32'h41f91a6a} /* (30, 23, 27) {real, imag} */,
  {32'hc198a3ef, 32'h42b598b9} /* (30, 23, 26) {real, imag} */,
  {32'hc19a3ba0, 32'hc2d43521} /* (30, 23, 25) {real, imag} */,
  {32'h4197a611, 32'h420314aa} /* (30, 23, 24) {real, imag} */,
  {32'h3f39bf50, 32'h4292acbe} /* (30, 23, 23) {real, imag} */,
  {32'hc09684d0, 32'hc28507fc} /* (30, 23, 22) {real, imag} */,
  {32'h40e6fe28, 32'h41e66186} /* (30, 23, 21) {real, imag} */,
  {32'hc22f1a2b, 32'hc0ab2040} /* (30, 23, 20) {real, imag} */,
  {32'h429374f0, 32'h4183dc0b} /* (30, 23, 19) {real, imag} */,
  {32'h420efb21, 32'h4265ed5c} /* (30, 23, 18) {real, imag} */,
  {32'h4277a1ca, 32'hc1b1bf7e} /* (30, 23, 17) {real, imag} */,
  {32'h41ba36f0, 32'h00000000} /* (30, 23, 16) {real, imag} */,
  {32'h4277a1ca, 32'h41b1bf7e} /* (30, 23, 15) {real, imag} */,
  {32'h420efb21, 32'hc265ed5c} /* (30, 23, 14) {real, imag} */,
  {32'h429374f0, 32'hc183dc0b} /* (30, 23, 13) {real, imag} */,
  {32'hc22f1a2b, 32'h40ab2040} /* (30, 23, 12) {real, imag} */,
  {32'h40e6fe28, 32'hc1e66186} /* (30, 23, 11) {real, imag} */,
  {32'hc09684d0, 32'h428507fc} /* (30, 23, 10) {real, imag} */,
  {32'h3f39bf50, 32'hc292acbe} /* (30, 23, 9) {real, imag} */,
  {32'h4197a611, 32'hc20314aa} /* (30, 23, 8) {real, imag} */,
  {32'hc19a3ba0, 32'h42d43521} /* (30, 23, 7) {real, imag} */,
  {32'hc198a3ef, 32'hc2b598b9} /* (30, 23, 6) {real, imag} */,
  {32'hc31a834e, 32'hc1f91a6a} /* (30, 23, 5) {real, imag} */,
  {32'h42d78c41, 32'h42e43a0a} /* (30, 23, 4) {real, imag} */,
  {32'h4318d446, 32'hc22536c8} /* (30, 23, 3) {real, imag} */,
  {32'hc4258a3f, 32'hc3a6be8b} /* (30, 23, 2) {real, imag} */,
  {32'h449257fa, 32'hc2866420} /* (30, 23, 1) {real, imag} */,
  {32'h44729179, 32'h00000000} /* (30, 23, 0) {real, imag} */,
  {32'h4446ca20, 32'h42c81025} /* (30, 22, 31) {real, imag} */,
  {32'hc4134e96, 32'h43b16e46} /* (30, 22, 30) {real, imag} */,
  {32'h433854ce, 32'h42c03046} /* (30, 22, 29) {real, imag} */,
  {32'hc19b4efc, 32'hc31104d4} /* (30, 22, 28) {real, imag} */,
  {32'hc344ba58, 32'h4037cdd0} /* (30, 22, 27) {real, imag} */,
  {32'hc262e9f4, 32'h41c61352} /* (30, 22, 26) {real, imag} */,
  {32'h42047f7a, 32'hc24cebb7} /* (30, 22, 25) {real, imag} */,
  {32'hc28cd7f6, 32'h428c944b} /* (30, 22, 24) {real, imag} */,
  {32'h41888ce0, 32'h42420f1a} /* (30, 22, 23) {real, imag} */,
  {32'h42898fbb, 32'h425145b8} /* (30, 22, 22) {real, imag} */,
  {32'hc28da602, 32'h42242264} /* (30, 22, 21) {real, imag} */,
  {32'hc23f633e, 32'hc01d9e00} /* (30, 22, 20) {real, imag} */,
  {32'h429ecb43, 32'hc22033f7} /* (30, 22, 19) {real, imag} */,
  {32'h426e5540, 32'hbfe4a260} /* (30, 22, 18) {real, imag} */,
  {32'hc2076580, 32'h3fe4daa0} /* (30, 22, 17) {real, imag} */,
  {32'h4212a3d5, 32'h00000000} /* (30, 22, 16) {real, imag} */,
  {32'hc2076580, 32'hbfe4daa0} /* (30, 22, 15) {real, imag} */,
  {32'h426e5540, 32'h3fe4a260} /* (30, 22, 14) {real, imag} */,
  {32'h429ecb43, 32'h422033f7} /* (30, 22, 13) {real, imag} */,
  {32'hc23f633e, 32'h401d9e00} /* (30, 22, 12) {real, imag} */,
  {32'hc28da602, 32'hc2242264} /* (30, 22, 11) {real, imag} */,
  {32'h42898fbb, 32'hc25145b8} /* (30, 22, 10) {real, imag} */,
  {32'h41888ce0, 32'hc2420f1a} /* (30, 22, 9) {real, imag} */,
  {32'hc28cd7f6, 32'hc28c944b} /* (30, 22, 8) {real, imag} */,
  {32'h42047f7a, 32'h424cebb7} /* (30, 22, 7) {real, imag} */,
  {32'hc262e9f4, 32'hc1c61352} /* (30, 22, 6) {real, imag} */,
  {32'hc344ba58, 32'hc037cdd0} /* (30, 22, 5) {real, imag} */,
  {32'hc19b4efc, 32'h431104d4} /* (30, 22, 4) {real, imag} */,
  {32'h433854ce, 32'hc2c03046} /* (30, 22, 3) {real, imag} */,
  {32'hc4134e96, 32'hc3b16e46} /* (30, 22, 2) {real, imag} */,
  {32'h4446ca20, 32'hc2c81025} /* (30, 22, 1) {real, imag} */,
  {32'h4426a97c, 32'h00000000} /* (30, 22, 0) {real, imag} */,
  {32'h432e56ca, 32'h434e35d1} /* (30, 21, 31) {real, imag} */,
  {32'hc3669951, 32'h42b00cc4} /* (30, 21, 30) {real, imag} */,
  {32'h42d10698, 32'h429dff73} /* (30, 21, 29) {real, imag} */,
  {32'hc1d4b9ee, 32'h42944c80} /* (30, 21, 28) {real, imag} */,
  {32'hc227463c, 32'hc1e2a9a5} /* (30, 21, 27) {real, imag} */,
  {32'hc2521d81, 32'hc275c02a} /* (30, 21, 26) {real, imag} */,
  {32'h42449380, 32'h41ad257a} /* (30, 21, 25) {real, imag} */,
  {32'hc2990c84, 32'hc16c46e8} /* (30, 21, 24) {real, imag} */,
  {32'hc192b018, 32'h417e8b2c} /* (30, 21, 23) {real, imag} */,
  {32'hbda80f00, 32'h422a8ad4} /* (30, 21, 22) {real, imag} */,
  {32'h42364742, 32'h41eef334} /* (30, 21, 21) {real, imag} */,
  {32'hc24b4b82, 32'h418fb3ef} /* (30, 21, 20) {real, imag} */,
  {32'hc2f8a22a, 32'h405a1a00} /* (30, 21, 19) {real, imag} */,
  {32'h4252bee4, 32'hc2751837} /* (30, 21, 18) {real, imag} */,
  {32'h424a352b, 32'h41625ae9} /* (30, 21, 17) {real, imag} */,
  {32'hc0db2428, 32'h00000000} /* (30, 21, 16) {real, imag} */,
  {32'h424a352b, 32'hc1625ae9} /* (30, 21, 15) {real, imag} */,
  {32'h4252bee4, 32'h42751837} /* (30, 21, 14) {real, imag} */,
  {32'hc2f8a22a, 32'hc05a1a00} /* (30, 21, 13) {real, imag} */,
  {32'hc24b4b82, 32'hc18fb3ef} /* (30, 21, 12) {real, imag} */,
  {32'h42364742, 32'hc1eef334} /* (30, 21, 11) {real, imag} */,
  {32'hbda80f00, 32'hc22a8ad4} /* (30, 21, 10) {real, imag} */,
  {32'hc192b018, 32'hc17e8b2c} /* (30, 21, 9) {real, imag} */,
  {32'hc2990c84, 32'h416c46e8} /* (30, 21, 8) {real, imag} */,
  {32'h42449380, 32'hc1ad257a} /* (30, 21, 7) {real, imag} */,
  {32'hc2521d81, 32'h4275c02a} /* (30, 21, 6) {real, imag} */,
  {32'hc227463c, 32'h41e2a9a5} /* (30, 21, 5) {real, imag} */,
  {32'hc1d4b9ee, 32'hc2944c80} /* (30, 21, 4) {real, imag} */,
  {32'h42d10698, 32'hc29dff73} /* (30, 21, 3) {real, imag} */,
  {32'hc3669951, 32'hc2b00cc4} /* (30, 21, 2) {real, imag} */,
  {32'h432e56ca, 32'hc34e35d1} /* (30, 21, 1) {real, imag} */,
  {32'h42823e70, 32'h00000000} /* (30, 21, 0) {real, imag} */,
  {32'hc45b8ec2, 32'h433d81c9} /* (30, 20, 31) {real, imag} */,
  {32'h43e7172a, 32'hc393b590} /* (30, 20, 30) {real, imag} */,
  {32'h4310c410, 32'h427a9154} /* (30, 20, 29) {real, imag} */,
  {32'hc31d33eb, 32'h425b51b6} /* (30, 20, 28) {real, imag} */,
  {32'h42a6cec2, 32'hc202f519} /* (30, 20, 27) {real, imag} */,
  {32'h421ce81b, 32'hc1bfb8c3} /* (30, 20, 26) {real, imag} */,
  {32'hc1adc952, 32'hc2067b42} /* (30, 20, 25) {real, imag} */,
  {32'hc2871bb2, 32'h42a62900} /* (30, 20, 24) {real, imag} */,
  {32'hc2cb6b12, 32'hc1b125e7} /* (30, 20, 23) {real, imag} */,
  {32'h412627fa, 32'hc245765c} /* (30, 20, 22) {real, imag} */,
  {32'hc20f2124, 32'hc2c723ff} /* (30, 20, 21) {real, imag} */,
  {32'hc2f54bba, 32'hc10f012a} /* (30, 20, 20) {real, imag} */,
  {32'h429d95eb, 32'h4280f269} /* (30, 20, 19) {real, imag} */,
  {32'h429697aa, 32'h41271274} /* (30, 20, 18) {real, imag} */,
  {32'h41c79dfa, 32'hc1904c04} /* (30, 20, 17) {real, imag} */,
  {32'hc2da65de, 32'h00000000} /* (30, 20, 16) {real, imag} */,
  {32'h41c79dfa, 32'h41904c04} /* (30, 20, 15) {real, imag} */,
  {32'h429697aa, 32'hc1271274} /* (30, 20, 14) {real, imag} */,
  {32'h429d95eb, 32'hc280f269} /* (30, 20, 13) {real, imag} */,
  {32'hc2f54bba, 32'h410f012a} /* (30, 20, 12) {real, imag} */,
  {32'hc20f2124, 32'h42c723ff} /* (30, 20, 11) {real, imag} */,
  {32'h412627fa, 32'h4245765c} /* (30, 20, 10) {real, imag} */,
  {32'hc2cb6b12, 32'h41b125e7} /* (30, 20, 9) {real, imag} */,
  {32'hc2871bb2, 32'hc2a62900} /* (30, 20, 8) {real, imag} */,
  {32'hc1adc952, 32'h42067b42} /* (30, 20, 7) {real, imag} */,
  {32'h421ce81b, 32'h41bfb8c3} /* (30, 20, 6) {real, imag} */,
  {32'h42a6cec2, 32'h4202f519} /* (30, 20, 5) {real, imag} */,
  {32'hc31d33eb, 32'hc25b51b6} /* (30, 20, 4) {real, imag} */,
  {32'h4310c410, 32'hc27a9154} /* (30, 20, 3) {real, imag} */,
  {32'h43e7172a, 32'h4393b590} /* (30, 20, 2) {real, imag} */,
  {32'hc45b8ec2, 32'hc33d81c9} /* (30, 20, 1) {real, imag} */,
  {32'hc43c40d6, 32'h00000000} /* (30, 20, 0) {real, imag} */,
  {32'hc4b31b67, 32'h42f9681a} /* (30, 19, 31) {real, imag} */,
  {32'h442e924b, 32'hc3b1721a} /* (30, 19, 30) {real, imag} */,
  {32'h42b14b02, 32'h42f3715b} /* (30, 19, 29) {real, imag} */,
  {32'hc3842553, 32'h42617159} /* (30, 19, 28) {real, imag} */,
  {32'h431746e8, 32'hc32cd7fc} /* (30, 19, 27) {real, imag} */,
  {32'h4270342c, 32'h418a834d} /* (30, 19, 26) {real, imag} */,
  {32'h411c50e8, 32'h41e38c24} /* (30, 19, 25) {real, imag} */,
  {32'hc21b1ed2, 32'hc245e8a8} /* (30, 19, 24) {real, imag} */,
  {32'h40f1291c, 32'h41db0bc9} /* (30, 19, 23) {real, imag} */,
  {32'hc2360614, 32'hc208daf1} /* (30, 19, 22) {real, imag} */,
  {32'hc15b34ec, 32'hc2f5ad48} /* (30, 19, 21) {real, imag} */,
  {32'h4028a460, 32'hc2bedf88} /* (30, 19, 20) {real, imag} */,
  {32'h42ca9bc0, 32'h420f5f9f} /* (30, 19, 19) {real, imag} */,
  {32'hc081a980, 32'hc22fa3d9} /* (30, 19, 18) {real, imag} */,
  {32'hc196d5eb, 32'h41c034f6} /* (30, 19, 17) {real, imag} */,
  {32'hc1e78ac3, 32'h00000000} /* (30, 19, 16) {real, imag} */,
  {32'hc196d5eb, 32'hc1c034f6} /* (30, 19, 15) {real, imag} */,
  {32'hc081a980, 32'h422fa3d9} /* (30, 19, 14) {real, imag} */,
  {32'h42ca9bc0, 32'hc20f5f9f} /* (30, 19, 13) {real, imag} */,
  {32'h4028a460, 32'h42bedf88} /* (30, 19, 12) {real, imag} */,
  {32'hc15b34ec, 32'h42f5ad48} /* (30, 19, 11) {real, imag} */,
  {32'hc2360614, 32'h4208daf1} /* (30, 19, 10) {real, imag} */,
  {32'h40f1291c, 32'hc1db0bc9} /* (30, 19, 9) {real, imag} */,
  {32'hc21b1ed2, 32'h4245e8a8} /* (30, 19, 8) {real, imag} */,
  {32'h411c50e8, 32'hc1e38c24} /* (30, 19, 7) {real, imag} */,
  {32'h4270342c, 32'hc18a834d} /* (30, 19, 6) {real, imag} */,
  {32'h431746e8, 32'h432cd7fc} /* (30, 19, 5) {real, imag} */,
  {32'hc3842553, 32'hc2617159} /* (30, 19, 4) {real, imag} */,
  {32'h42b14b02, 32'hc2f3715b} /* (30, 19, 3) {real, imag} */,
  {32'h442e924b, 32'h43b1721a} /* (30, 19, 2) {real, imag} */,
  {32'hc4b31b67, 32'hc2f9681a} /* (30, 19, 1) {real, imag} */,
  {32'hc47f735e, 32'h00000000} /* (30, 19, 0) {real, imag} */,
  {32'hc4cd0918, 32'hc1c611a0} /* (30, 18, 31) {real, imag} */,
  {32'h44268f4d, 32'hc35fc4aa} /* (30, 18, 30) {real, imag} */,
  {32'h4216b73b, 32'h436a85d3} /* (30, 18, 29) {real, imag} */,
  {32'hc3877c7e, 32'h42a44c72} /* (30, 18, 28) {real, imag} */,
  {32'h434b0ac5, 32'hc36e463b} /* (30, 18, 27) {real, imag} */,
  {32'h412ae650, 32'h42f3c866} /* (30, 18, 26) {real, imag} */,
  {32'hc208bdf4, 32'h42de1a0d} /* (30, 18, 25) {real, imag} */,
  {32'h4270c3cf, 32'hc07acf40} /* (30, 18, 24) {real, imag} */,
  {32'h422d25ec, 32'h428ecc4e} /* (30, 18, 23) {real, imag} */,
  {32'hc2180838, 32'hc1c1008e} /* (30, 18, 22) {real, imag} */,
  {32'h4290ae03, 32'hc2dd60fc} /* (30, 18, 21) {real, imag} */,
  {32'h427eba70, 32'h428e2a33} /* (30, 18, 20) {real, imag} */,
  {32'hc213f78c, 32'h41168f78} /* (30, 18, 19) {real, imag} */,
  {32'h40480a1c, 32'hc19d3f72} /* (30, 18, 18) {real, imag} */,
  {32'h4265283f, 32'hc21704a5} /* (30, 18, 17) {real, imag} */,
  {32'h4125dbb8, 32'h00000000} /* (30, 18, 16) {real, imag} */,
  {32'h4265283f, 32'h421704a5} /* (30, 18, 15) {real, imag} */,
  {32'h40480a1c, 32'h419d3f72} /* (30, 18, 14) {real, imag} */,
  {32'hc213f78c, 32'hc1168f78} /* (30, 18, 13) {real, imag} */,
  {32'h427eba70, 32'hc28e2a33} /* (30, 18, 12) {real, imag} */,
  {32'h4290ae03, 32'h42dd60fc} /* (30, 18, 11) {real, imag} */,
  {32'hc2180838, 32'h41c1008e} /* (30, 18, 10) {real, imag} */,
  {32'h422d25ec, 32'hc28ecc4e} /* (30, 18, 9) {real, imag} */,
  {32'h4270c3cf, 32'h407acf40} /* (30, 18, 8) {real, imag} */,
  {32'hc208bdf4, 32'hc2de1a0d} /* (30, 18, 7) {real, imag} */,
  {32'h412ae650, 32'hc2f3c866} /* (30, 18, 6) {real, imag} */,
  {32'h434b0ac5, 32'h436e463b} /* (30, 18, 5) {real, imag} */,
  {32'hc3877c7e, 32'hc2a44c72} /* (30, 18, 4) {real, imag} */,
  {32'h4216b73b, 32'hc36a85d3} /* (30, 18, 3) {real, imag} */,
  {32'h44268f4d, 32'h435fc4aa} /* (30, 18, 2) {real, imag} */,
  {32'hc4cd0918, 32'h41c611a0} /* (30, 18, 1) {real, imag} */,
  {32'hc4869ff3, 32'h00000000} /* (30, 18, 0) {real, imag} */,
  {32'hc4de3232, 32'h4221dad4} /* (30, 17, 31) {real, imag} */,
  {32'h442433f7, 32'hc341182a} /* (30, 17, 30) {real, imag} */,
  {32'h408c49d8, 32'h43207550} /* (30, 17, 29) {real, imag} */,
  {32'hc32397fc, 32'h42e3aa31} /* (30, 17, 28) {real, imag} */,
  {32'h435c3fb8, 32'hc2f3dda5} /* (30, 17, 27) {real, imag} */,
  {32'h3fcf94e0, 32'h428c4e9f} /* (30, 17, 26) {real, imag} */,
  {32'hc299e7a2, 32'h4275cc54} /* (30, 17, 25) {real, imag} */,
  {32'h424bcbf9, 32'hc23513dc} /* (30, 17, 24) {real, imag} */,
  {32'h421f263e, 32'h41ed9a66} /* (30, 17, 23) {real, imag} */,
  {32'hbf1b74a0, 32'h42cdcc3e} /* (30, 17, 22) {real, imag} */,
  {32'h42c417fa, 32'hc32881f3} /* (30, 17, 21) {real, imag} */,
  {32'hc12f1092, 32'h414e033e} /* (30, 17, 20) {real, imag} */,
  {32'hc1b26fd3, 32'hc0bb3920} /* (30, 17, 19) {real, imag} */,
  {32'h41bef18a, 32'hc246ec59} /* (30, 17, 18) {real, imag} */,
  {32'h3dc09300, 32'h42c20126} /* (30, 17, 17) {real, imag} */,
  {32'hc1eeb35a, 32'h00000000} /* (30, 17, 16) {real, imag} */,
  {32'h3dc09300, 32'hc2c20126} /* (30, 17, 15) {real, imag} */,
  {32'h41bef18a, 32'h4246ec59} /* (30, 17, 14) {real, imag} */,
  {32'hc1b26fd3, 32'h40bb3920} /* (30, 17, 13) {real, imag} */,
  {32'hc12f1092, 32'hc14e033e} /* (30, 17, 12) {real, imag} */,
  {32'h42c417fa, 32'h432881f3} /* (30, 17, 11) {real, imag} */,
  {32'hbf1b74a0, 32'hc2cdcc3e} /* (30, 17, 10) {real, imag} */,
  {32'h421f263e, 32'hc1ed9a66} /* (30, 17, 9) {real, imag} */,
  {32'h424bcbf9, 32'h423513dc} /* (30, 17, 8) {real, imag} */,
  {32'hc299e7a2, 32'hc275cc54} /* (30, 17, 7) {real, imag} */,
  {32'h3fcf94e0, 32'hc28c4e9f} /* (30, 17, 6) {real, imag} */,
  {32'h435c3fb8, 32'h42f3dda5} /* (30, 17, 5) {real, imag} */,
  {32'hc32397fc, 32'hc2e3aa31} /* (30, 17, 4) {real, imag} */,
  {32'h408c49d8, 32'hc3207550} /* (30, 17, 3) {real, imag} */,
  {32'h442433f7, 32'h4341182a} /* (30, 17, 2) {real, imag} */,
  {32'hc4de3232, 32'hc221dad4} /* (30, 17, 1) {real, imag} */,
  {32'hc4914448, 32'h00000000} /* (30, 17, 0) {real, imag} */,
  {32'hc4e254ff, 32'hc18e7540} /* (30, 16, 31) {real, imag} */,
  {32'h444ccf9c, 32'hc2f2b916} /* (30, 16, 30) {real, imag} */,
  {32'hc10c0844, 32'hc281b163} /* (30, 16, 29) {real, imag} */,
  {32'hc3494726, 32'h428a0240} /* (30, 16, 28) {real, imag} */,
  {32'h43873877, 32'h42eb9e58} /* (30, 16, 27) {real, imag} */,
  {32'h42570dda, 32'h419297bc} /* (30, 16, 26) {real, imag} */,
  {32'hc17d8658, 32'hc2cb0bfd} /* (30, 16, 25) {real, imag} */,
  {32'h43072472, 32'hc2c9bdef} /* (30, 16, 24) {real, imag} */,
  {32'hbeff6c40, 32'h42d83773} /* (30, 16, 23) {real, imag} */,
  {32'h41569112, 32'hc2740ec6} /* (30, 16, 22) {real, imag} */,
  {32'hc044ba20, 32'hc2c995f4} /* (30, 16, 21) {real, imag} */,
  {32'hc2a13814, 32'h4237f743} /* (30, 16, 20) {real, imag} */,
  {32'h412a80c2, 32'h4288b2c6} /* (30, 16, 19) {real, imag} */,
  {32'h427434be, 32'h42070e62} /* (30, 16, 18) {real, imag} */,
  {32'h424467a0, 32'hc25b38bd} /* (30, 16, 17) {real, imag} */,
  {32'hc292c86a, 32'h00000000} /* (30, 16, 16) {real, imag} */,
  {32'h424467a0, 32'h425b38bd} /* (30, 16, 15) {real, imag} */,
  {32'h427434be, 32'hc2070e62} /* (30, 16, 14) {real, imag} */,
  {32'h412a80c2, 32'hc288b2c6} /* (30, 16, 13) {real, imag} */,
  {32'hc2a13814, 32'hc237f743} /* (30, 16, 12) {real, imag} */,
  {32'hc044ba20, 32'h42c995f4} /* (30, 16, 11) {real, imag} */,
  {32'h41569112, 32'h42740ec6} /* (30, 16, 10) {real, imag} */,
  {32'hbeff6c40, 32'hc2d83773} /* (30, 16, 9) {real, imag} */,
  {32'h43072472, 32'h42c9bdef} /* (30, 16, 8) {real, imag} */,
  {32'hc17d8658, 32'h42cb0bfd} /* (30, 16, 7) {real, imag} */,
  {32'h42570dda, 32'hc19297bc} /* (30, 16, 6) {real, imag} */,
  {32'h43873877, 32'hc2eb9e58} /* (30, 16, 5) {real, imag} */,
  {32'hc3494726, 32'hc28a0240} /* (30, 16, 4) {real, imag} */,
  {32'hc10c0844, 32'h4281b163} /* (30, 16, 3) {real, imag} */,
  {32'h444ccf9c, 32'h42f2b916} /* (30, 16, 2) {real, imag} */,
  {32'hc4e254ff, 32'h418e7540} /* (30, 16, 1) {real, imag} */,
  {32'hc4a148ab, 32'h00000000} /* (30, 16, 0) {real, imag} */,
  {32'hc4d0c1a2, 32'hc2dcfd22} /* (30, 15, 31) {real, imag} */,
  {32'h44544331, 32'hc3063d7a} /* (30, 15, 30) {real, imag} */,
  {32'hc1e0cf0a, 32'h42d71a41} /* (30, 15, 29) {real, imag} */,
  {32'hc242198c, 32'h425e731a} /* (30, 15, 28) {real, imag} */,
  {32'h43503f00, 32'h40d93890} /* (30, 15, 27) {real, imag} */,
  {32'h408a6f08, 32'h3ffd2a40} /* (30, 15, 26) {real, imag} */,
  {32'h412f26e0, 32'hc14fcda0} /* (30, 15, 25) {real, imag} */,
  {32'hc1ba756a, 32'hc3030193} /* (30, 15, 24) {real, imag} */,
  {32'h4160a901, 32'h4164d3b5} /* (30, 15, 23) {real, imag} */,
  {32'h4218caca, 32'hc0ffa408} /* (30, 15, 22) {real, imag} */,
  {32'h41f128f8, 32'h41ff5178} /* (30, 15, 21) {real, imag} */,
  {32'h41b8c23f, 32'hc1b91a2d} /* (30, 15, 20) {real, imag} */,
  {32'hc2a186a3, 32'hc259294d} /* (30, 15, 19) {real, imag} */,
  {32'h41883cee, 32'hc0f1dc08} /* (30, 15, 18) {real, imag} */,
  {32'h4267543c, 32'hc1eb5a26} /* (30, 15, 17) {real, imag} */,
  {32'h412eba05, 32'h00000000} /* (30, 15, 16) {real, imag} */,
  {32'h4267543c, 32'h41eb5a26} /* (30, 15, 15) {real, imag} */,
  {32'h41883cee, 32'h40f1dc08} /* (30, 15, 14) {real, imag} */,
  {32'hc2a186a3, 32'h4259294d} /* (30, 15, 13) {real, imag} */,
  {32'h41b8c23f, 32'h41b91a2d} /* (30, 15, 12) {real, imag} */,
  {32'h41f128f8, 32'hc1ff5178} /* (30, 15, 11) {real, imag} */,
  {32'h4218caca, 32'h40ffa408} /* (30, 15, 10) {real, imag} */,
  {32'h4160a901, 32'hc164d3b5} /* (30, 15, 9) {real, imag} */,
  {32'hc1ba756a, 32'h43030193} /* (30, 15, 8) {real, imag} */,
  {32'h412f26e0, 32'h414fcda0} /* (30, 15, 7) {real, imag} */,
  {32'h408a6f08, 32'hbffd2a40} /* (30, 15, 6) {real, imag} */,
  {32'h43503f00, 32'hc0d93890} /* (30, 15, 5) {real, imag} */,
  {32'hc242198c, 32'hc25e731a} /* (30, 15, 4) {real, imag} */,
  {32'hc1e0cf0a, 32'hc2d71a41} /* (30, 15, 3) {real, imag} */,
  {32'h44544331, 32'h43063d7a} /* (30, 15, 2) {real, imag} */,
  {32'hc4d0c1a2, 32'h42dcfd22} /* (30, 15, 1) {real, imag} */,
  {32'hc4a9d3b8, 32'h00000000} /* (30, 15, 0) {real, imag} */,
  {32'hc4bba010, 32'hc1aaf020} /* (30, 14, 31) {real, imag} */,
  {32'h4453babb, 32'hc303b202} /* (30, 14, 30) {real, imag} */,
  {32'hc13aa3bc, 32'h43081961} /* (30, 14, 29) {real, imag} */,
  {32'hc2d47eba, 32'h42c62e52} /* (30, 14, 28) {real, imag} */,
  {32'h432bf0d7, 32'h427b5194} /* (30, 14, 27) {real, imag} */,
  {32'h42eccb4c, 32'h41fab60a} /* (30, 14, 26) {real, imag} */,
  {32'hc1bdf1ef, 32'h42b7334b} /* (30, 14, 25) {real, imag} */,
  {32'h41e5ba52, 32'hc2e920fe} /* (30, 14, 24) {real, imag} */,
  {32'h4151d3cf, 32'hc0d50e08} /* (30, 14, 23) {real, imag} */,
  {32'h41a48ace, 32'h427d8c2f} /* (30, 14, 22) {real, imag} */,
  {32'h42192e5a, 32'h421c1d67} /* (30, 14, 21) {real, imag} */,
  {32'hc146be46, 32'hc23429aa} /* (30, 14, 20) {real, imag} */,
  {32'hc289ecba, 32'h425cf488} /* (30, 14, 19) {real, imag} */,
  {32'hc11f43e9, 32'hc2d36a26} /* (30, 14, 18) {real, imag} */,
  {32'hc242763d, 32'h41d4fe6e} /* (30, 14, 17) {real, imag} */,
  {32'h420aa920, 32'h00000000} /* (30, 14, 16) {real, imag} */,
  {32'hc242763d, 32'hc1d4fe6e} /* (30, 14, 15) {real, imag} */,
  {32'hc11f43e9, 32'h42d36a26} /* (30, 14, 14) {real, imag} */,
  {32'hc289ecba, 32'hc25cf488} /* (30, 14, 13) {real, imag} */,
  {32'hc146be46, 32'h423429aa} /* (30, 14, 12) {real, imag} */,
  {32'h42192e5a, 32'hc21c1d67} /* (30, 14, 11) {real, imag} */,
  {32'h41a48ace, 32'hc27d8c2f} /* (30, 14, 10) {real, imag} */,
  {32'h4151d3cf, 32'h40d50e08} /* (30, 14, 9) {real, imag} */,
  {32'h41e5ba52, 32'h42e920fe} /* (30, 14, 8) {real, imag} */,
  {32'hc1bdf1ef, 32'hc2b7334b} /* (30, 14, 7) {real, imag} */,
  {32'h42eccb4c, 32'hc1fab60a} /* (30, 14, 6) {real, imag} */,
  {32'h432bf0d7, 32'hc27b5194} /* (30, 14, 5) {real, imag} */,
  {32'hc2d47eba, 32'hc2c62e52} /* (30, 14, 4) {real, imag} */,
  {32'hc13aa3bc, 32'hc3081961} /* (30, 14, 3) {real, imag} */,
  {32'h4453babb, 32'h4303b202} /* (30, 14, 2) {real, imag} */,
  {32'hc4bba010, 32'h41aaf020} /* (30, 14, 1) {real, imag} */,
  {32'hc4a2b867, 32'h00000000} /* (30, 14, 0) {real, imag} */,
  {32'hc4b040bb, 32'h41ce2ab8} /* (30, 13, 31) {real, imag} */,
  {32'h445e455d, 32'hc33efae4} /* (30, 13, 30) {real, imag} */,
  {32'h420e74b0, 32'hc1b09a94} /* (30, 13, 29) {real, imag} */,
  {32'hc2be7c3c, 32'h430b8a06} /* (30, 13, 28) {real, imag} */,
  {32'h42d5e4c4, 32'h4287e3b4} /* (30, 13, 27) {real, imag} */,
  {32'h429d38a0, 32'hc17e29c6} /* (30, 13, 26) {real, imag} */,
  {32'hc30ccef0, 32'h42d35107} /* (30, 13, 25) {real, imag} */,
  {32'hc1fd540d, 32'hc22b8c38} /* (30, 13, 24) {real, imag} */,
  {32'h412fd3a2, 32'h422e3798} /* (30, 13, 23) {real, imag} */,
  {32'h424d4efc, 32'hc15d43e4} /* (30, 13, 22) {real, imag} */,
  {32'hc0aabf48, 32'hc2faa8ae} /* (30, 13, 21) {real, imag} */,
  {32'hc2a78ccf, 32'h41ad35e2} /* (30, 13, 20) {real, imag} */,
  {32'h4226c3e0, 32'hc240877d} /* (30, 13, 19) {real, imag} */,
  {32'hc18b8a16, 32'hc285cfba} /* (30, 13, 18) {real, imag} */,
  {32'h42222560, 32'hbf0d3830} /* (30, 13, 17) {real, imag} */,
  {32'h420a1228, 32'h00000000} /* (30, 13, 16) {real, imag} */,
  {32'h42222560, 32'h3f0d3830} /* (30, 13, 15) {real, imag} */,
  {32'hc18b8a16, 32'h4285cfba} /* (30, 13, 14) {real, imag} */,
  {32'h4226c3e0, 32'h4240877d} /* (30, 13, 13) {real, imag} */,
  {32'hc2a78ccf, 32'hc1ad35e2} /* (30, 13, 12) {real, imag} */,
  {32'hc0aabf48, 32'h42faa8ae} /* (30, 13, 11) {real, imag} */,
  {32'h424d4efc, 32'h415d43e4} /* (30, 13, 10) {real, imag} */,
  {32'h412fd3a2, 32'hc22e3798} /* (30, 13, 9) {real, imag} */,
  {32'hc1fd540d, 32'h422b8c38} /* (30, 13, 8) {real, imag} */,
  {32'hc30ccef0, 32'hc2d35107} /* (30, 13, 7) {real, imag} */,
  {32'h429d38a0, 32'h417e29c6} /* (30, 13, 6) {real, imag} */,
  {32'h42d5e4c4, 32'hc287e3b4} /* (30, 13, 5) {real, imag} */,
  {32'hc2be7c3c, 32'hc30b8a06} /* (30, 13, 4) {real, imag} */,
  {32'h420e74b0, 32'h41b09a94} /* (30, 13, 3) {real, imag} */,
  {32'h445e455d, 32'h433efae4} /* (30, 13, 2) {real, imag} */,
  {32'hc4b040bb, 32'hc1ce2ab8} /* (30, 13, 1) {real, imag} */,
  {32'hc4b2da65, 32'h00000000} /* (30, 13, 0) {real, imag} */,
  {32'hc49007fc, 32'h4272f724} /* (30, 12, 31) {real, imag} */,
  {32'h443038e9, 32'hc33a6e8b} /* (30, 12, 30) {real, imag} */,
  {32'hc1fa88cc, 32'hc2d23992} /* (30, 12, 29) {real, imag} */,
  {32'hc25f65cc, 32'h4279197e} /* (30, 12, 28) {real, imag} */,
  {32'h42e7b8aa, 32'hc2e4eeb0} /* (30, 12, 27) {real, imag} */,
  {32'hc2933aca, 32'h422c4636} /* (30, 12, 26) {real, imag} */,
  {32'hc15bd544, 32'h42b74c74} /* (30, 12, 25) {real, imag} */,
  {32'h41a811a2, 32'h41001750} /* (30, 12, 24) {real, imag} */,
  {32'hc26b122d, 32'h42079886} /* (30, 12, 23) {real, imag} */,
  {32'hc0c5aac4, 32'hc15e92d0} /* (30, 12, 22) {real, imag} */,
  {32'hc18b5040, 32'hc20ec64a} /* (30, 12, 21) {real, imag} */,
  {32'hc1cd8fb6, 32'hc22a1f44} /* (30, 12, 20) {real, imag} */,
  {32'hc2297776, 32'h4189ac7d} /* (30, 12, 19) {real, imag} */,
  {32'hc186c0ff, 32'h422363a9} /* (30, 12, 18) {real, imag} */,
  {32'h4173b488, 32'h419b02e6} /* (30, 12, 17) {real, imag} */,
  {32'hc148e56c, 32'h00000000} /* (30, 12, 16) {real, imag} */,
  {32'h4173b488, 32'hc19b02e6} /* (30, 12, 15) {real, imag} */,
  {32'hc186c0ff, 32'hc22363a9} /* (30, 12, 14) {real, imag} */,
  {32'hc2297776, 32'hc189ac7d} /* (30, 12, 13) {real, imag} */,
  {32'hc1cd8fb6, 32'h422a1f44} /* (30, 12, 12) {real, imag} */,
  {32'hc18b5040, 32'h420ec64a} /* (30, 12, 11) {real, imag} */,
  {32'hc0c5aac4, 32'h415e92d0} /* (30, 12, 10) {real, imag} */,
  {32'hc26b122d, 32'hc2079886} /* (30, 12, 9) {real, imag} */,
  {32'h41a811a2, 32'hc1001750} /* (30, 12, 8) {real, imag} */,
  {32'hc15bd544, 32'hc2b74c74} /* (30, 12, 7) {real, imag} */,
  {32'hc2933aca, 32'hc22c4636} /* (30, 12, 6) {real, imag} */,
  {32'h42e7b8aa, 32'h42e4eeb0} /* (30, 12, 5) {real, imag} */,
  {32'hc25f65cc, 32'hc279197e} /* (30, 12, 4) {real, imag} */,
  {32'hc1fa88cc, 32'h42d23992} /* (30, 12, 3) {real, imag} */,
  {32'h443038e9, 32'h433a6e8b} /* (30, 12, 2) {real, imag} */,
  {32'hc49007fc, 32'hc272f724} /* (30, 12, 1) {real, imag} */,
  {32'hc49092ab, 32'h00000000} /* (30, 12, 0) {real, imag} */,
  {32'hc429331c, 32'h42644dbc} /* (30, 11, 31) {real, imag} */,
  {32'h43fcb6ee, 32'hc1b218e0} /* (30, 11, 30) {real, imag} */,
  {32'hc3034400, 32'hc237f904} /* (30, 11, 29) {real, imag} */,
  {32'hc0fd8798, 32'hc1f70113} /* (30, 11, 28) {real, imag} */,
  {32'h42fa1728, 32'hc2abd694} /* (30, 11, 27) {real, imag} */,
  {32'h425a4779, 32'h414abe08} /* (30, 11, 26) {real, imag} */,
  {32'hc228e22a, 32'h4290a042} /* (30, 11, 25) {real, imag} */,
  {32'h41d3ba32, 32'hc2fd453d} /* (30, 11, 24) {real, imag} */,
  {32'hc2a2fd7e, 32'hc1fe092e} /* (30, 11, 23) {real, imag} */,
  {32'hc25bb13a, 32'h43715ff7} /* (30, 11, 22) {real, imag} */,
  {32'hc274aa0e, 32'hc20421fc} /* (30, 11, 21) {real, imag} */,
  {32'h4254217a, 32'hc27a34d0} /* (30, 11, 20) {real, imag} */,
  {32'hc2bb4aae, 32'hc2ab3d68} /* (30, 11, 19) {real, imag} */,
  {32'h41436dce, 32'h41cc4e9e} /* (30, 11, 18) {real, imag} */,
  {32'h423f1791, 32'hc1c42174} /* (30, 11, 17) {real, imag} */,
  {32'h423e19b7, 32'h00000000} /* (30, 11, 16) {real, imag} */,
  {32'h423f1791, 32'h41c42174} /* (30, 11, 15) {real, imag} */,
  {32'h41436dce, 32'hc1cc4e9e} /* (30, 11, 14) {real, imag} */,
  {32'hc2bb4aae, 32'h42ab3d68} /* (30, 11, 13) {real, imag} */,
  {32'h4254217a, 32'h427a34d0} /* (30, 11, 12) {real, imag} */,
  {32'hc274aa0e, 32'h420421fc} /* (30, 11, 11) {real, imag} */,
  {32'hc25bb13a, 32'hc3715ff7} /* (30, 11, 10) {real, imag} */,
  {32'hc2a2fd7e, 32'h41fe092e} /* (30, 11, 9) {real, imag} */,
  {32'h41d3ba32, 32'h42fd453d} /* (30, 11, 8) {real, imag} */,
  {32'hc228e22a, 32'hc290a042} /* (30, 11, 7) {real, imag} */,
  {32'h425a4779, 32'hc14abe08} /* (30, 11, 6) {real, imag} */,
  {32'h42fa1728, 32'h42abd694} /* (30, 11, 5) {real, imag} */,
  {32'hc0fd8798, 32'h41f70113} /* (30, 11, 4) {real, imag} */,
  {32'hc3034400, 32'h4237f904} /* (30, 11, 3) {real, imag} */,
  {32'h43fcb6ee, 32'h41b218e0} /* (30, 11, 2) {real, imag} */,
  {32'hc429331c, 32'hc2644dbc} /* (30, 11, 1) {real, imag} */,
  {32'hc41504f0, 32'h00000000} /* (30, 11, 0) {real, imag} */,
  {32'h43e51c20, 32'h4210120e} /* (30, 10, 31) {real, imag} */,
  {32'hc3288678, 32'h43527f03} /* (30, 10, 30) {real, imag} */,
  {32'hc2c2b0f0, 32'hc2949fb6} /* (30, 10, 29) {real, imag} */,
  {32'h42faf1d1, 32'hc188936e} /* (30, 10, 28) {real, imag} */,
  {32'h40c761b0, 32'hc2d87ee8} /* (30, 10, 27) {real, imag} */,
  {32'h4203ec6e, 32'hbf4d3ab0} /* (30, 10, 26) {real, imag} */,
  {32'hc21a4d82, 32'hc2193ef1} /* (30, 10, 25) {real, imag} */,
  {32'hc283f08e, 32'hc2cda19d} /* (30, 10, 24) {real, imag} */,
  {32'h41ea0932, 32'h41a09cc4} /* (30, 10, 23) {real, imag} */,
  {32'h40ec47f0, 32'h4287632c} /* (30, 10, 22) {real, imag} */,
  {32'hc1f36eb4, 32'hc1c83b48} /* (30, 10, 21) {real, imag} */,
  {32'hc28fd4d8, 32'h4290ef90} /* (30, 10, 20) {real, imag} */,
  {32'hc1dc0ceb, 32'h40ee8bb0} /* (30, 10, 19) {real, imag} */,
  {32'hc0f41880, 32'hc275841b} /* (30, 10, 18) {real, imag} */,
  {32'h41340076, 32'hc23e9c3a} /* (30, 10, 17) {real, imag} */,
  {32'h4233c78d, 32'h00000000} /* (30, 10, 16) {real, imag} */,
  {32'h41340076, 32'h423e9c3a} /* (30, 10, 15) {real, imag} */,
  {32'hc0f41880, 32'h4275841b} /* (30, 10, 14) {real, imag} */,
  {32'hc1dc0ceb, 32'hc0ee8bb0} /* (30, 10, 13) {real, imag} */,
  {32'hc28fd4d8, 32'hc290ef90} /* (30, 10, 12) {real, imag} */,
  {32'hc1f36eb4, 32'h41c83b48} /* (30, 10, 11) {real, imag} */,
  {32'h40ec47f0, 32'hc287632c} /* (30, 10, 10) {real, imag} */,
  {32'h41ea0932, 32'hc1a09cc4} /* (30, 10, 9) {real, imag} */,
  {32'hc283f08e, 32'h42cda19d} /* (30, 10, 8) {real, imag} */,
  {32'hc21a4d82, 32'h42193ef1} /* (30, 10, 7) {real, imag} */,
  {32'h4203ec6e, 32'h3f4d3ab0} /* (30, 10, 6) {real, imag} */,
  {32'h40c761b0, 32'h42d87ee8} /* (30, 10, 5) {real, imag} */,
  {32'h42faf1d1, 32'h4188936e} /* (30, 10, 4) {real, imag} */,
  {32'hc2c2b0f0, 32'h42949fb6} /* (30, 10, 3) {real, imag} */,
  {32'hc3288678, 32'hc3527f03} /* (30, 10, 2) {real, imag} */,
  {32'h43e51c20, 32'hc210120e} /* (30, 10, 1) {real, imag} */,
  {32'h434559e5, 32'h00000000} /* (30, 10, 0) {real, imag} */,
  {32'h4494f304, 32'hc2e6d254} /* (30, 9, 31) {real, imag} */,
  {32'hc3d314ae, 32'h43847efd} /* (30, 9, 30) {real, imag} */,
  {32'hc165ff80, 32'hc01ecc78} /* (30, 9, 29) {real, imag} */,
  {32'h420641c6, 32'hc10e7c44} /* (30, 9, 28) {real, imag} */,
  {32'hc1a13700, 32'h4191323a} /* (30, 9, 27) {real, imag} */,
  {32'hc220d4f6, 32'hc118dc20} /* (30, 9, 26) {real, imag} */,
  {32'h41d72900, 32'hc15efc68} /* (30, 9, 25) {real, imag} */,
  {32'hc276422c, 32'h42b50f40} /* (30, 9, 24) {real, imag} */,
  {32'h40c02f4e, 32'h41ec043e} /* (30, 9, 23) {real, imag} */,
  {32'hc2ac8037, 32'hc1bbddce} /* (30, 9, 22) {real, imag} */,
  {32'hc1965ace, 32'h428d9cdc} /* (30, 9, 21) {real, imag} */,
  {32'hc1684ccc, 32'hc2150709} /* (30, 9, 20) {real, imag} */,
  {32'h42b9991c, 32'h42841c23} /* (30, 9, 19) {real, imag} */,
  {32'h420fa6b5, 32'h42a32e1e} /* (30, 9, 18) {real, imag} */,
  {32'h41222836, 32'h4278ee35} /* (30, 9, 17) {real, imag} */,
  {32'hc2b99dc2, 32'h00000000} /* (30, 9, 16) {real, imag} */,
  {32'h41222836, 32'hc278ee35} /* (30, 9, 15) {real, imag} */,
  {32'h420fa6b5, 32'hc2a32e1e} /* (30, 9, 14) {real, imag} */,
  {32'h42b9991c, 32'hc2841c23} /* (30, 9, 13) {real, imag} */,
  {32'hc1684ccc, 32'h42150709} /* (30, 9, 12) {real, imag} */,
  {32'hc1965ace, 32'hc28d9cdc} /* (30, 9, 11) {real, imag} */,
  {32'hc2ac8037, 32'h41bbddce} /* (30, 9, 10) {real, imag} */,
  {32'h40c02f4e, 32'hc1ec043e} /* (30, 9, 9) {real, imag} */,
  {32'hc276422c, 32'hc2b50f40} /* (30, 9, 8) {real, imag} */,
  {32'h41d72900, 32'h415efc68} /* (30, 9, 7) {real, imag} */,
  {32'hc220d4f6, 32'h4118dc20} /* (30, 9, 6) {real, imag} */,
  {32'hc1a13700, 32'hc191323a} /* (30, 9, 5) {real, imag} */,
  {32'h420641c6, 32'h410e7c44} /* (30, 9, 4) {real, imag} */,
  {32'hc165ff80, 32'h401ecc78} /* (30, 9, 3) {real, imag} */,
  {32'hc3d314ae, 32'hc3847efd} /* (30, 9, 2) {real, imag} */,
  {32'h4494f304, 32'h42e6d254} /* (30, 9, 1) {real, imag} */,
  {32'h44075467, 32'h00000000} /* (30, 9, 0) {real, imag} */,
  {32'h44c2193a, 32'hc39356a4} /* (30, 8, 31) {real, imag} */,
  {32'hc401b462, 32'h43bcf034} /* (30, 8, 30) {real, imag} */,
  {32'hc294dac4, 32'hc1c194bb} /* (30, 8, 29) {real, imag} */,
  {32'h4308962b, 32'h41d9d550} /* (30, 8, 28) {real, imag} */,
  {32'hc32ce2be, 32'h4289e1e6} /* (30, 8, 27) {real, imag} */,
  {32'h4031aca0, 32'hc24d9325} /* (30, 8, 26) {real, imag} */,
  {32'hc1cde51c, 32'hc1b85bb0} /* (30, 8, 25) {real, imag} */,
  {32'hc2e4cdaa, 32'h41f2cb46} /* (30, 8, 24) {real, imag} */,
  {32'h4164ccac, 32'hc1bf0610} /* (30, 8, 23) {real, imag} */,
  {32'h42c9b2e9, 32'h41065f4c} /* (30, 8, 22) {real, imag} */,
  {32'hbfae5500, 32'h42d1700c} /* (30, 8, 21) {real, imag} */,
  {32'h42b2cbce, 32'hc20d68d6} /* (30, 8, 20) {real, imag} */,
  {32'hc219a16a, 32'h423f74cd} /* (30, 8, 19) {real, imag} */,
  {32'hc218f81f, 32'hc20ba321} /* (30, 8, 18) {real, imag} */,
  {32'h429afaa8, 32'h426f1da1} /* (30, 8, 17) {real, imag} */,
  {32'hc2fb0862, 32'h00000000} /* (30, 8, 16) {real, imag} */,
  {32'h429afaa8, 32'hc26f1da1} /* (30, 8, 15) {real, imag} */,
  {32'hc218f81f, 32'h420ba321} /* (30, 8, 14) {real, imag} */,
  {32'hc219a16a, 32'hc23f74cd} /* (30, 8, 13) {real, imag} */,
  {32'h42b2cbce, 32'h420d68d6} /* (30, 8, 12) {real, imag} */,
  {32'hbfae5500, 32'hc2d1700c} /* (30, 8, 11) {real, imag} */,
  {32'h42c9b2e9, 32'hc1065f4c} /* (30, 8, 10) {real, imag} */,
  {32'h4164ccac, 32'h41bf0610} /* (30, 8, 9) {real, imag} */,
  {32'hc2e4cdaa, 32'hc1f2cb46} /* (30, 8, 8) {real, imag} */,
  {32'hc1cde51c, 32'h41b85bb0} /* (30, 8, 7) {real, imag} */,
  {32'h4031aca0, 32'h424d9325} /* (30, 8, 6) {real, imag} */,
  {32'hc32ce2be, 32'hc289e1e6} /* (30, 8, 5) {real, imag} */,
  {32'h4308962b, 32'hc1d9d550} /* (30, 8, 4) {real, imag} */,
  {32'hc294dac4, 32'h41c194bb} /* (30, 8, 3) {real, imag} */,
  {32'hc401b462, 32'hc3bcf034} /* (30, 8, 2) {real, imag} */,
  {32'h44c2193a, 32'h439356a4} /* (30, 8, 1) {real, imag} */,
  {32'h43e53d7c, 32'h00000000} /* (30, 8, 0) {real, imag} */,
  {32'h44bf7809, 32'hc3360d46} /* (30, 7, 31) {real, imag} */,
  {32'hc3f58014, 32'h43eed588} /* (30, 7, 30) {real, imag} */,
  {32'hc2fb48c0, 32'h42883798} /* (30, 7, 29) {real, imag} */,
  {32'h43252b70, 32'hc1c2f151} /* (30, 7, 28) {real, imag} */,
  {32'hc31940c5, 32'h429afd42} /* (30, 7, 27) {real, imag} */,
  {32'hc238ea92, 32'h40a059b0} /* (30, 7, 26) {real, imag} */,
  {32'h42a9c6bb, 32'hc03d40c0} /* (30, 7, 25) {real, imag} */,
  {32'hc29863ba, 32'h41cece57} /* (30, 7, 24) {real, imag} */,
  {32'hc0cbcebe, 32'hc234137f} /* (30, 7, 23) {real, imag} */,
  {32'h4242ca34, 32'hc2bdd154} /* (30, 7, 22) {real, imag} */,
  {32'hc2c7025e, 32'hc1fa519c} /* (30, 7, 21) {real, imag} */,
  {32'hc242aed8, 32'hc22c110a} /* (30, 7, 20) {real, imag} */,
  {32'h421c2488, 32'h40000438} /* (30, 7, 19) {real, imag} */,
  {32'hc20bd38f, 32'h423b2b25} /* (30, 7, 18) {real, imag} */,
  {32'hc058e758, 32'h408c01da} /* (30, 7, 17) {real, imag} */,
  {32'hc11c7ed6, 32'h00000000} /* (30, 7, 16) {real, imag} */,
  {32'hc058e758, 32'hc08c01da} /* (30, 7, 15) {real, imag} */,
  {32'hc20bd38f, 32'hc23b2b25} /* (30, 7, 14) {real, imag} */,
  {32'h421c2488, 32'hc0000438} /* (30, 7, 13) {real, imag} */,
  {32'hc242aed8, 32'h422c110a} /* (30, 7, 12) {real, imag} */,
  {32'hc2c7025e, 32'h41fa519c} /* (30, 7, 11) {real, imag} */,
  {32'h4242ca34, 32'h42bdd154} /* (30, 7, 10) {real, imag} */,
  {32'hc0cbcebe, 32'h4234137f} /* (30, 7, 9) {real, imag} */,
  {32'hc29863ba, 32'hc1cece57} /* (30, 7, 8) {real, imag} */,
  {32'h42a9c6bb, 32'h403d40c0} /* (30, 7, 7) {real, imag} */,
  {32'hc238ea92, 32'hc0a059b0} /* (30, 7, 6) {real, imag} */,
  {32'hc31940c5, 32'hc29afd42} /* (30, 7, 5) {real, imag} */,
  {32'h43252b70, 32'h41c2f151} /* (30, 7, 4) {real, imag} */,
  {32'hc2fb48c0, 32'hc2883798} /* (30, 7, 3) {real, imag} */,
  {32'hc3f58014, 32'hc3eed588} /* (30, 7, 2) {real, imag} */,
  {32'h44bf7809, 32'h43360d46} /* (30, 7, 1) {real, imag} */,
  {32'h444361e0, 32'h00000000} /* (30, 7, 0) {real, imag} */,
  {32'h44a76a60, 32'hc3b795fe} /* (30, 6, 31) {real, imag} */,
  {32'hc3f1750c, 32'h43faa71e} /* (30, 6, 30) {real, imag} */,
  {32'h41ffc7e6, 32'h3e053d00} /* (30, 6, 29) {real, imag} */,
  {32'h4319be17, 32'hc2caec8c} /* (30, 6, 28) {real, imag} */,
  {32'hc2e1595c, 32'h428698ed} /* (30, 6, 27) {real, imag} */,
  {32'hc318fd6a, 32'h42650ab8} /* (30, 6, 26) {real, imag} */,
  {32'hc16610e2, 32'h421693d0} /* (30, 6, 25) {real, imag} */,
  {32'hc2078665, 32'h42e7fde8} /* (30, 6, 24) {real, imag} */,
  {32'hc286e432, 32'hc2136cca} /* (30, 6, 23) {real, imag} */,
  {32'h42804654, 32'hc30e0eba} /* (30, 6, 22) {real, imag} */,
  {32'hc1e4f97e, 32'h4319e462} /* (30, 6, 21) {real, imag} */,
  {32'h413dd90c, 32'hc2a71d06} /* (30, 6, 20) {real, imag} */,
  {32'h4213ffe2, 32'hc1aa4a71} /* (30, 6, 19) {real, imag} */,
  {32'h421eba80, 32'hc21f054b} /* (30, 6, 18) {real, imag} */,
  {32'h40b82864, 32'h413aea26} /* (30, 6, 17) {real, imag} */,
  {32'hc2bc0852, 32'h00000000} /* (30, 6, 16) {real, imag} */,
  {32'h40b82864, 32'hc13aea26} /* (30, 6, 15) {real, imag} */,
  {32'h421eba80, 32'h421f054b} /* (30, 6, 14) {real, imag} */,
  {32'h4213ffe2, 32'h41aa4a71} /* (30, 6, 13) {real, imag} */,
  {32'h413dd90c, 32'h42a71d06} /* (30, 6, 12) {real, imag} */,
  {32'hc1e4f97e, 32'hc319e462} /* (30, 6, 11) {real, imag} */,
  {32'h42804654, 32'h430e0eba} /* (30, 6, 10) {real, imag} */,
  {32'hc286e432, 32'h42136cca} /* (30, 6, 9) {real, imag} */,
  {32'hc2078665, 32'hc2e7fde8} /* (30, 6, 8) {real, imag} */,
  {32'hc16610e2, 32'hc21693d0} /* (30, 6, 7) {real, imag} */,
  {32'hc318fd6a, 32'hc2650ab8} /* (30, 6, 6) {real, imag} */,
  {32'hc2e1595c, 32'hc28698ed} /* (30, 6, 5) {real, imag} */,
  {32'h4319be17, 32'h42caec8c} /* (30, 6, 4) {real, imag} */,
  {32'h41ffc7e6, 32'hbe053d00} /* (30, 6, 3) {real, imag} */,
  {32'hc3f1750c, 32'hc3faa71e} /* (30, 6, 2) {real, imag} */,
  {32'h44a76a60, 32'h43b795fe} /* (30, 6, 1) {real, imag} */,
  {32'h44381878, 32'h00000000} /* (30, 6, 0) {real, imag} */,
  {32'h4488925e, 32'hc44a9406} /* (30, 5, 31) {real, imag} */,
  {32'hc2f35854, 32'h44210e35} /* (30, 5, 30) {real, imag} */,
  {32'hc2078cab, 32'hc1856ab8} /* (30, 5, 29) {real, imag} */,
  {32'hc28720ba, 32'h41bd2f76} /* (30, 5, 28) {real, imag} */,
  {32'hc30208e2, 32'h416e88be} /* (30, 5, 27) {real, imag} */,
  {32'hc2859582, 32'hc1a3ba7c} /* (30, 5, 26) {real, imag} */,
  {32'h41754640, 32'h423a37bb} /* (30, 5, 25) {real, imag} */,
  {32'h4276a770, 32'h42ddb486} /* (30, 5, 24) {real, imag} */,
  {32'hc24c383d, 32'hc109a484} /* (30, 5, 23) {real, imag} */,
  {32'h41a0f2cd, 32'h40d1a368} /* (30, 5, 22) {real, imag} */,
  {32'hc1c1d797, 32'hc1ec668a} /* (30, 5, 21) {real, imag} */,
  {32'hbe81dc80, 32'hc24ce0f2} /* (30, 5, 20) {real, imag} */,
  {32'hc2836052, 32'hc1a26390} /* (30, 5, 19) {real, imag} */,
  {32'h410c363a, 32'h41856cd2} /* (30, 5, 18) {real, imag} */,
  {32'h4146e86a, 32'h427f898b} /* (30, 5, 17) {real, imag} */,
  {32'h42c24ae2, 32'h00000000} /* (30, 5, 16) {real, imag} */,
  {32'h4146e86a, 32'hc27f898b} /* (30, 5, 15) {real, imag} */,
  {32'h410c363a, 32'hc1856cd2} /* (30, 5, 14) {real, imag} */,
  {32'hc2836052, 32'h41a26390} /* (30, 5, 13) {real, imag} */,
  {32'hbe81dc80, 32'h424ce0f2} /* (30, 5, 12) {real, imag} */,
  {32'hc1c1d797, 32'h41ec668a} /* (30, 5, 11) {real, imag} */,
  {32'h41a0f2cd, 32'hc0d1a368} /* (30, 5, 10) {real, imag} */,
  {32'hc24c383d, 32'h4109a484} /* (30, 5, 9) {real, imag} */,
  {32'h4276a770, 32'hc2ddb486} /* (30, 5, 8) {real, imag} */,
  {32'h41754640, 32'hc23a37bb} /* (30, 5, 7) {real, imag} */,
  {32'hc2859582, 32'h41a3ba7c} /* (30, 5, 6) {real, imag} */,
  {32'hc30208e2, 32'hc16e88be} /* (30, 5, 5) {real, imag} */,
  {32'hc28720ba, 32'hc1bd2f76} /* (30, 5, 4) {real, imag} */,
  {32'hc2078cab, 32'h41856ab8} /* (30, 5, 3) {real, imag} */,
  {32'hc2f35854, 32'hc4210e35} /* (30, 5, 2) {real, imag} */,
  {32'h4488925e, 32'h444a9406} /* (30, 5, 1) {real, imag} */,
  {32'h4434f976, 32'h00000000} /* (30, 5, 0) {real, imag} */,
  {32'h44452738, 32'hc4877ed6} /* (30, 4, 31) {real, imag} */,
  {32'h42b44fe8, 32'h443c3232} /* (30, 4, 30) {real, imag} */,
  {32'hc35716bc, 32'hc002ec50} /* (30, 4, 29) {real, imag} */,
  {32'hc323ec40, 32'h41e38bdb} /* (30, 4, 28) {real, imag} */,
  {32'hc19b97d0, 32'h421e941e} /* (30, 4, 27) {real, imag} */,
  {32'hbfca26f0, 32'h4230b574} /* (30, 4, 26) {real, imag} */,
  {32'h40ca32d8, 32'hc25aad3c} /* (30, 4, 25) {real, imag} */,
  {32'h42aba8ff, 32'h41556e78} /* (30, 4, 24) {real, imag} */,
  {32'hc0987f1a, 32'hc18ad09a} /* (30, 4, 23) {real, imag} */,
  {32'h41f6ecd2, 32'hc09e047e} /* (30, 4, 22) {real, imag} */,
  {32'hc10af0fc, 32'hc21b7564} /* (30, 4, 21) {real, imag} */,
  {32'h42059c7f, 32'h424c551c} /* (30, 4, 20) {real, imag} */,
  {32'hc18bdac1, 32'h4201ae46} /* (30, 4, 19) {real, imag} */,
  {32'h425ddc7a, 32'h42c5851c} /* (30, 4, 18) {real, imag} */,
  {32'hc2605db7, 32'h423ea624} /* (30, 4, 17) {real, imag} */,
  {32'h4010a8f0, 32'h00000000} /* (30, 4, 16) {real, imag} */,
  {32'hc2605db7, 32'hc23ea624} /* (30, 4, 15) {real, imag} */,
  {32'h425ddc7a, 32'hc2c5851c} /* (30, 4, 14) {real, imag} */,
  {32'hc18bdac1, 32'hc201ae46} /* (30, 4, 13) {real, imag} */,
  {32'h42059c7f, 32'hc24c551c} /* (30, 4, 12) {real, imag} */,
  {32'hc10af0fc, 32'h421b7564} /* (30, 4, 11) {real, imag} */,
  {32'h41f6ecd2, 32'h409e047e} /* (30, 4, 10) {real, imag} */,
  {32'hc0987f1a, 32'h418ad09a} /* (30, 4, 9) {real, imag} */,
  {32'h42aba8ff, 32'hc1556e78} /* (30, 4, 8) {real, imag} */,
  {32'h40ca32d8, 32'h425aad3c} /* (30, 4, 7) {real, imag} */,
  {32'hbfca26f0, 32'hc230b574} /* (30, 4, 6) {real, imag} */,
  {32'hc19b97d0, 32'hc21e941e} /* (30, 4, 5) {real, imag} */,
  {32'hc323ec40, 32'hc1e38bdb} /* (30, 4, 4) {real, imag} */,
  {32'hc35716bc, 32'h4002ec50} /* (30, 4, 3) {real, imag} */,
  {32'h42b44fe8, 32'hc43c3232} /* (30, 4, 2) {real, imag} */,
  {32'h44452738, 32'h44877ed6} /* (30, 4, 1) {real, imag} */,
  {32'h44189924, 32'h00000000} /* (30, 4, 0) {real, imag} */,
  {32'h443a6dbb, 32'hc4a5d0ec} /* (30, 3, 31) {real, imag} */,
  {32'h432d18e4, 32'h442931a8} /* (30, 3, 30) {real, imag} */,
  {32'hc28907d6, 32'h42310f36} /* (30, 3, 29) {real, imag} */,
  {32'hc29269a5, 32'h43055439} /* (30, 3, 28) {real, imag} */,
  {32'hc2fa0e86, 32'h42e62f06} /* (30, 3, 27) {real, imag} */,
  {32'hc1a9eb20, 32'hc2bb33c2} /* (30, 3, 26) {real, imag} */,
  {32'hc211f527, 32'hc3084cb0} /* (30, 3, 25) {real, imag} */,
  {32'hc2bbf523, 32'h43471738} /* (30, 3, 24) {real, imag} */,
  {32'hc2339005, 32'hc2044964} /* (30, 3, 23) {real, imag} */,
  {32'hc1285b8a, 32'h428ae64f} /* (30, 3, 22) {real, imag} */,
  {32'hc25b8a75, 32'hc1f976fc} /* (30, 3, 21) {real, imag} */,
  {32'h42896842, 32'hc19593b2} /* (30, 3, 20) {real, imag} */,
  {32'hc1c7f34b, 32'hc2452b35} /* (30, 3, 19) {real, imag} */,
  {32'hc1b90ac9, 32'hc30f9538} /* (30, 3, 18) {real, imag} */,
  {32'h42890a11, 32'h40dddde0} /* (30, 3, 17) {real, imag} */,
  {32'hc16b246c, 32'h00000000} /* (30, 3, 16) {real, imag} */,
  {32'h42890a11, 32'hc0dddde0} /* (30, 3, 15) {real, imag} */,
  {32'hc1b90ac9, 32'h430f9538} /* (30, 3, 14) {real, imag} */,
  {32'hc1c7f34b, 32'h42452b35} /* (30, 3, 13) {real, imag} */,
  {32'h42896842, 32'h419593b2} /* (30, 3, 12) {real, imag} */,
  {32'hc25b8a75, 32'h41f976fc} /* (30, 3, 11) {real, imag} */,
  {32'hc1285b8a, 32'hc28ae64f} /* (30, 3, 10) {real, imag} */,
  {32'hc2339005, 32'h42044964} /* (30, 3, 9) {real, imag} */,
  {32'hc2bbf523, 32'hc3471738} /* (30, 3, 8) {real, imag} */,
  {32'hc211f527, 32'h43084cb0} /* (30, 3, 7) {real, imag} */,
  {32'hc1a9eb20, 32'h42bb33c2} /* (30, 3, 6) {real, imag} */,
  {32'hc2fa0e86, 32'hc2e62f06} /* (30, 3, 5) {real, imag} */,
  {32'hc29269a5, 32'hc3055439} /* (30, 3, 4) {real, imag} */,
  {32'hc28907d6, 32'hc2310f36} /* (30, 3, 3) {real, imag} */,
  {32'h432d18e4, 32'hc42931a8} /* (30, 3, 2) {real, imag} */,
  {32'h443a6dbb, 32'h44a5d0ec} /* (30, 3, 1) {real, imag} */,
  {32'h43fc264c, 32'h00000000} /* (30, 3, 0) {real, imag} */,
  {32'h441d0e60, 32'hc4a6db96} /* (30, 2, 31) {real, imag} */,
  {32'h4348c590, 32'h43f97a35} /* (30, 2, 30) {real, imag} */,
  {32'hc267f341, 32'h420c1358} /* (30, 2, 29) {real, imag} */,
  {32'hc32a5966, 32'h4313965e} /* (30, 2, 28) {real, imag} */,
  {32'hc2e3f9a0, 32'h41caf3b8} /* (30, 2, 27) {real, imag} */,
  {32'hc2c2d0ce, 32'hc2b58c7e} /* (30, 2, 26) {real, imag} */,
  {32'hc1aa141d, 32'hc2c968b5} /* (30, 2, 25) {real, imag} */,
  {32'h41e418f6, 32'h42f168f4} /* (30, 2, 24) {real, imag} */,
  {32'hc18e9cca, 32'hc0d0ed58} /* (30, 2, 23) {real, imag} */,
  {32'hc1030286, 32'h42b2ee22} /* (30, 2, 22) {real, imag} */,
  {32'hc01eda00, 32'hc25bacfc} /* (30, 2, 21) {real, imag} */,
  {32'h429bcd6e, 32'hc221b156} /* (30, 2, 20) {real, imag} */,
  {32'hc291e7c7, 32'h41715302} /* (30, 2, 19) {real, imag} */,
  {32'hc26493e2, 32'h42aaa72c} /* (30, 2, 18) {real, imag} */,
  {32'h4224f242, 32'h420e39ca} /* (30, 2, 17) {real, imag} */,
  {32'h427c6fa4, 32'h00000000} /* (30, 2, 16) {real, imag} */,
  {32'h4224f242, 32'hc20e39ca} /* (30, 2, 15) {real, imag} */,
  {32'hc26493e2, 32'hc2aaa72c} /* (30, 2, 14) {real, imag} */,
  {32'hc291e7c7, 32'hc1715302} /* (30, 2, 13) {real, imag} */,
  {32'h429bcd6e, 32'h4221b156} /* (30, 2, 12) {real, imag} */,
  {32'hc01eda00, 32'h425bacfc} /* (30, 2, 11) {real, imag} */,
  {32'hc1030286, 32'hc2b2ee22} /* (30, 2, 10) {real, imag} */,
  {32'hc18e9cca, 32'h40d0ed58} /* (30, 2, 9) {real, imag} */,
  {32'h41e418f6, 32'hc2f168f4} /* (30, 2, 8) {real, imag} */,
  {32'hc1aa141d, 32'h42c968b5} /* (30, 2, 7) {real, imag} */,
  {32'hc2c2d0ce, 32'h42b58c7e} /* (30, 2, 6) {real, imag} */,
  {32'hc2e3f9a0, 32'hc1caf3b8} /* (30, 2, 5) {real, imag} */,
  {32'hc32a5966, 32'hc313965e} /* (30, 2, 4) {real, imag} */,
  {32'hc267f341, 32'hc20c1358} /* (30, 2, 3) {real, imag} */,
  {32'h4348c590, 32'hc3f97a35} /* (30, 2, 2) {real, imag} */,
  {32'h441d0e60, 32'h44a6db96} /* (30, 2, 1) {real, imag} */,
  {32'h439d9804, 32'h00000000} /* (30, 2, 0) {real, imag} */,
  {32'h44001c50, 32'hc491b9c6} /* (30, 1, 31) {real, imag} */,
  {32'h4314636c, 32'h440bff6c} /* (30, 1, 30) {real, imag} */,
  {32'hc2b034ec, 32'h4224e5c8} /* (30, 1, 29) {real, imag} */,
  {32'hc2c9c6b5, 32'h43253b3a} /* (30, 1, 28) {real, imag} */,
  {32'hc2c0e6d1, 32'hc285eb4a} /* (30, 1, 27) {real, imag} */,
  {32'hc2f6fedc, 32'hbf167220} /* (30, 1, 26) {real, imag} */,
  {32'hc1d1642c, 32'hc33a2a4a} /* (30, 1, 25) {real, imag} */,
  {32'h4152b638, 32'h42eeaafd} /* (30, 1, 24) {real, imag} */,
  {32'h424e903f, 32'hc20481ad} /* (30, 1, 23) {real, imag} */,
  {32'h416ddae2, 32'h41a6d681} /* (30, 1, 22) {real, imag} */,
  {32'hc2ac3bd4, 32'h414cdd64} /* (30, 1, 21) {real, imag} */,
  {32'hc0e32cf9, 32'h42577852} /* (30, 1, 20) {real, imag} */,
  {32'h42b7920c, 32'hc2ee1a55} /* (30, 1, 19) {real, imag} */,
  {32'h41ac354e, 32'h425ce5a1} /* (30, 1, 18) {real, imag} */,
  {32'hc0e386ac, 32'hc14d98b4} /* (30, 1, 17) {real, imag} */,
  {32'hc1fc61b8, 32'h00000000} /* (30, 1, 16) {real, imag} */,
  {32'hc0e386ac, 32'h414d98b4} /* (30, 1, 15) {real, imag} */,
  {32'h41ac354e, 32'hc25ce5a1} /* (30, 1, 14) {real, imag} */,
  {32'h42b7920c, 32'h42ee1a55} /* (30, 1, 13) {real, imag} */,
  {32'hc0e32cf9, 32'hc2577852} /* (30, 1, 12) {real, imag} */,
  {32'hc2ac3bd4, 32'hc14cdd64} /* (30, 1, 11) {real, imag} */,
  {32'h416ddae2, 32'hc1a6d681} /* (30, 1, 10) {real, imag} */,
  {32'h424e903f, 32'h420481ad} /* (30, 1, 9) {real, imag} */,
  {32'h4152b638, 32'hc2eeaafd} /* (30, 1, 8) {real, imag} */,
  {32'hc1d1642c, 32'h433a2a4a} /* (30, 1, 7) {real, imag} */,
  {32'hc2f6fedc, 32'h3f167220} /* (30, 1, 6) {real, imag} */,
  {32'hc2c0e6d1, 32'h4285eb4a} /* (30, 1, 5) {real, imag} */,
  {32'hc2c9c6b5, 32'hc3253b3a} /* (30, 1, 4) {real, imag} */,
  {32'hc2b034ec, 32'hc224e5c8} /* (30, 1, 3) {real, imag} */,
  {32'h4314636c, 32'hc40bff6c} /* (30, 1, 2) {real, imag} */,
  {32'h44001c50, 32'h4491b9c6} /* (30, 1, 1) {real, imag} */,
  {32'h43b16c62, 32'h00000000} /* (30, 1, 0) {real, imag} */,
  {32'h4407ae0e, 32'hc457a7da} /* (30, 0, 31) {real, imag} */,
  {32'hc2de05a0, 32'h43fe4f10} /* (30, 0, 30) {real, imag} */,
  {32'hc1fe739c, 32'hc180562c} /* (30, 0, 29) {real, imag} */,
  {32'hc17d9ae8, 32'h43345ee7} /* (30, 0, 28) {real, imag} */,
  {32'hc30eb8b3, 32'hc2ab2fbe} /* (30, 0, 27) {real, imag} */,
  {32'h4284fc83, 32'hc1a1c94e} /* (30, 0, 26) {real, imag} */,
  {32'hc14114c8, 32'hc2cdb9bb} /* (30, 0, 25) {real, imag} */,
  {32'h40297ba0, 32'h423182de} /* (30, 0, 24) {real, imag} */,
  {32'hc05ff2a8, 32'hc0959cb0} /* (30, 0, 23) {real, imag} */,
  {32'hc1691bce, 32'hc2870e43} /* (30, 0, 22) {real, imag} */,
  {32'h402bef40, 32'h40054fb0} /* (30, 0, 21) {real, imag} */,
  {32'hc23a1ffb, 32'h41baefc2} /* (30, 0, 20) {real, imag} */,
  {32'hc1304c3e, 32'hc14f82cc} /* (30, 0, 19) {real, imag} */,
  {32'hc23e6790, 32'h41b096e1} /* (30, 0, 18) {real, imag} */,
  {32'h41b4ea84, 32'hc0c25290} /* (30, 0, 17) {real, imag} */,
  {32'h4116074c, 32'h00000000} /* (30, 0, 16) {real, imag} */,
  {32'h41b4ea84, 32'h40c25290} /* (30, 0, 15) {real, imag} */,
  {32'hc23e6790, 32'hc1b096e1} /* (30, 0, 14) {real, imag} */,
  {32'hc1304c3e, 32'h414f82cc} /* (30, 0, 13) {real, imag} */,
  {32'hc23a1ffb, 32'hc1baefc2} /* (30, 0, 12) {real, imag} */,
  {32'h402bef40, 32'hc0054fb0} /* (30, 0, 11) {real, imag} */,
  {32'hc1691bce, 32'h42870e43} /* (30, 0, 10) {real, imag} */,
  {32'hc05ff2a8, 32'h40959cb0} /* (30, 0, 9) {real, imag} */,
  {32'h40297ba0, 32'hc23182de} /* (30, 0, 8) {real, imag} */,
  {32'hc14114c8, 32'h42cdb9bb} /* (30, 0, 7) {real, imag} */,
  {32'h4284fc83, 32'h41a1c94e} /* (30, 0, 6) {real, imag} */,
  {32'hc30eb8b3, 32'h42ab2fbe} /* (30, 0, 5) {real, imag} */,
  {32'hc17d9ae8, 32'hc3345ee7} /* (30, 0, 4) {real, imag} */,
  {32'hc1fe739c, 32'h4180562c} /* (30, 0, 3) {real, imag} */,
  {32'hc2de05a0, 32'hc3fe4f10} /* (30, 0, 2) {real, imag} */,
  {32'h4407ae0e, 32'h4457a7da} /* (30, 0, 1) {real, imag} */,
  {32'h43b4e2a8, 32'h00000000} /* (30, 0, 0) {real, imag} */,
  {32'h44633da2, 32'hc40edabb} /* (29, 31, 31) {real, imag} */,
  {32'hc3dda059, 32'h43fcd1bd} /* (29, 31, 30) {real, imag} */,
  {32'hc21f1187, 32'hc248b96c} /* (29, 31, 29) {real, imag} */,
  {32'h42ce8922, 32'h42983d1f} /* (29, 31, 28) {real, imag} */,
  {32'hc302820f, 32'h42727082} /* (29, 31, 27) {real, imag} */,
  {32'hc23e845c, 32'hc15c906e} /* (29, 31, 26) {real, imag} */,
  {32'h41c4cdff, 32'h421239f4} /* (29, 31, 25) {real, imag} */,
  {32'hc1539930, 32'h4217e41a} /* (29, 31, 24) {real, imag} */,
  {32'hc1533b11, 32'hc0b7ef30} /* (29, 31, 23) {real, imag} */,
  {32'h428e89b6, 32'h4133bf8e} /* (29, 31, 22) {real, imag} */,
  {32'h41922c0a, 32'h4232f2f3} /* (29, 31, 21) {real, imag} */,
  {32'h3ff0ec38, 32'h4189d654} /* (29, 31, 20) {real, imag} */,
  {32'hc0e06ed4, 32'hc2849464} /* (29, 31, 19) {real, imag} */,
  {32'hc27d6f68, 32'hc20aa69b} /* (29, 31, 18) {real, imag} */,
  {32'h41995092, 32'h42298370} /* (29, 31, 17) {real, imag} */,
  {32'hc1cbbe10, 32'h00000000} /* (29, 31, 16) {real, imag} */,
  {32'h41995092, 32'hc2298370} /* (29, 31, 15) {real, imag} */,
  {32'hc27d6f68, 32'h420aa69b} /* (29, 31, 14) {real, imag} */,
  {32'hc0e06ed4, 32'h42849464} /* (29, 31, 13) {real, imag} */,
  {32'h3ff0ec38, 32'hc189d654} /* (29, 31, 12) {real, imag} */,
  {32'h41922c0a, 32'hc232f2f3} /* (29, 31, 11) {real, imag} */,
  {32'h428e89b6, 32'hc133bf8e} /* (29, 31, 10) {real, imag} */,
  {32'hc1533b11, 32'h40b7ef30} /* (29, 31, 9) {real, imag} */,
  {32'hc1539930, 32'hc217e41a} /* (29, 31, 8) {real, imag} */,
  {32'h41c4cdff, 32'hc21239f4} /* (29, 31, 7) {real, imag} */,
  {32'hc23e845c, 32'h415c906e} /* (29, 31, 6) {real, imag} */,
  {32'hc302820f, 32'hc2727082} /* (29, 31, 5) {real, imag} */,
  {32'h42ce8922, 32'hc2983d1f} /* (29, 31, 4) {real, imag} */,
  {32'hc21f1187, 32'h4248b96c} /* (29, 31, 3) {real, imag} */,
  {32'hc3dda059, 32'hc3fcd1bd} /* (29, 31, 2) {real, imag} */,
  {32'h44633da2, 32'h440edabb} /* (29, 31, 1) {real, imag} */,
  {32'h43d1a884, 32'h00000000} /* (29, 31, 0) {real, imag} */,
  {32'h44b3033e, 32'hc3db3d88} /* (29, 30, 31) {real, imag} */,
  {32'hc44c31f6, 32'h43f868eb} /* (29, 30, 30) {real, imag} */,
  {32'hc28609cd, 32'hc1022a70} /* (29, 30, 29) {real, imag} */,
  {32'h432d71d0, 32'h42ebc1de} /* (29, 30, 28) {real, imag} */,
  {32'hc3301171, 32'h432a965e} /* (29, 30, 27) {real, imag} */,
  {32'hc280d100, 32'hc214cc8c} /* (29, 30, 26) {real, imag} */,
  {32'h42758a93, 32'h41b7dcb0} /* (29, 30, 25) {real, imag} */,
  {32'h4106d10a, 32'h42c25920} /* (29, 30, 24) {real, imag} */,
  {32'hc13979e4, 32'h41e18d41} /* (29, 30, 23) {real, imag} */,
  {32'h428d78e7, 32'hc2af453f} /* (29, 30, 22) {real, imag} */,
  {32'h42903195, 32'h42a01d23} /* (29, 30, 21) {real, imag} */,
  {32'h40f1cc70, 32'h42eca77b} /* (29, 30, 20) {real, imag} */,
  {32'hc2160790, 32'h42a3006c} /* (29, 30, 19) {real, imag} */,
  {32'h41fc7e2c, 32'h40eaa073} /* (29, 30, 18) {real, imag} */,
  {32'h413ae68e, 32'hc20609ba} /* (29, 30, 17) {real, imag} */,
  {32'hc2339573, 32'h00000000} /* (29, 30, 16) {real, imag} */,
  {32'h413ae68e, 32'h420609ba} /* (29, 30, 15) {real, imag} */,
  {32'h41fc7e2c, 32'hc0eaa073} /* (29, 30, 14) {real, imag} */,
  {32'hc2160790, 32'hc2a3006c} /* (29, 30, 13) {real, imag} */,
  {32'h40f1cc70, 32'hc2eca77b} /* (29, 30, 12) {real, imag} */,
  {32'h42903195, 32'hc2a01d23} /* (29, 30, 11) {real, imag} */,
  {32'h428d78e7, 32'h42af453f} /* (29, 30, 10) {real, imag} */,
  {32'hc13979e4, 32'hc1e18d41} /* (29, 30, 9) {real, imag} */,
  {32'h4106d10a, 32'hc2c25920} /* (29, 30, 8) {real, imag} */,
  {32'h42758a93, 32'hc1b7dcb0} /* (29, 30, 7) {real, imag} */,
  {32'hc280d100, 32'h4214cc8c} /* (29, 30, 6) {real, imag} */,
  {32'hc3301171, 32'hc32a965e} /* (29, 30, 5) {real, imag} */,
  {32'h432d71d0, 32'hc2ebc1de} /* (29, 30, 4) {real, imag} */,
  {32'hc28609cd, 32'h41022a70} /* (29, 30, 3) {real, imag} */,
  {32'hc44c31f6, 32'hc3f868eb} /* (29, 30, 2) {real, imag} */,
  {32'h44b3033e, 32'h43db3d88} /* (29, 30, 1) {real, imag} */,
  {32'h44369d61, 32'h00000000} /* (29, 30, 0) {real, imag} */,
  {32'h44d4ee18, 32'hc3891154} /* (29, 29, 31) {real, imag} */,
  {32'hc4895838, 32'h43ae5637} /* (29, 29, 30) {real, imag} */,
  {32'h40799620, 32'hc282f6b3} /* (29, 29, 29) {real, imag} */,
  {32'h4378fd13, 32'h4240fd9c} /* (29, 29, 28) {real, imag} */,
  {32'hc363610a, 32'hc2f15cbd} /* (29, 29, 27) {real, imag} */,
  {32'h421a293c, 32'hc2a2bcc0} /* (29, 29, 26) {real, imag} */,
  {32'hc1c3e5a6, 32'hc27de5d6} /* (29, 29, 25) {real, imag} */,
  {32'hc12644de, 32'hc2df3221} /* (29, 29, 24) {real, imag} */,
  {32'hc2aeb6d8, 32'h42a323bf} /* (29, 29, 23) {real, imag} */,
  {32'hc0e503e0, 32'hc304aeaf} /* (29, 29, 22) {real, imag} */,
  {32'hc2052712, 32'h42dea344} /* (29, 29, 21) {real, imag} */,
  {32'h4255115c, 32'hc2188eae} /* (29, 29, 20) {real, imag} */,
  {32'hc3045b94, 32'h4264c46e} /* (29, 29, 19) {real, imag} */,
  {32'hc174c3d6, 32'h42c7260c} /* (29, 29, 18) {real, imag} */,
  {32'h421b30ac, 32'hc2905be5} /* (29, 29, 17) {real, imag} */,
  {32'hc2ba6b90, 32'h00000000} /* (29, 29, 16) {real, imag} */,
  {32'h421b30ac, 32'h42905be5} /* (29, 29, 15) {real, imag} */,
  {32'hc174c3d6, 32'hc2c7260c} /* (29, 29, 14) {real, imag} */,
  {32'hc3045b94, 32'hc264c46e} /* (29, 29, 13) {real, imag} */,
  {32'h4255115c, 32'h42188eae} /* (29, 29, 12) {real, imag} */,
  {32'hc2052712, 32'hc2dea344} /* (29, 29, 11) {real, imag} */,
  {32'hc0e503e0, 32'h4304aeaf} /* (29, 29, 10) {real, imag} */,
  {32'hc2aeb6d8, 32'hc2a323bf} /* (29, 29, 9) {real, imag} */,
  {32'hc12644de, 32'h42df3221} /* (29, 29, 8) {real, imag} */,
  {32'hc1c3e5a6, 32'h427de5d6} /* (29, 29, 7) {real, imag} */,
  {32'h421a293c, 32'h42a2bcc0} /* (29, 29, 6) {real, imag} */,
  {32'hc363610a, 32'h42f15cbd} /* (29, 29, 5) {real, imag} */,
  {32'h4378fd13, 32'hc240fd9c} /* (29, 29, 4) {real, imag} */,
  {32'h40799620, 32'h4282f6b3} /* (29, 29, 3) {real, imag} */,
  {32'hc4895838, 32'hc3ae5637} /* (29, 29, 2) {real, imag} */,
  {32'h44d4ee18, 32'h43891154} /* (29, 29, 1) {real, imag} */,
  {32'h441d77a4, 32'h00000000} /* (29, 29, 0) {real, imag} */,
  {32'h44cae112, 32'hc2c14650} /* (29, 28, 31) {real, imag} */,
  {32'hc48c409c, 32'h439a1c8c} /* (29, 28, 30) {real, imag} */,
  {32'hc0acd4a8, 32'hc3834130} /* (29, 28, 29) {real, imag} */,
  {32'h43593aca, 32'hc249ae6c} /* (29, 28, 28) {real, imag} */,
  {32'hc34b8a56, 32'h42d915de} /* (29, 28, 27) {real, imag} */,
  {32'h423b1904, 32'hc28315fb} /* (29, 28, 26) {real, imag} */,
  {32'hc2ce4658, 32'hc28dde02} /* (29, 28, 25) {real, imag} */,
  {32'hc09a5af0, 32'h423d77fc} /* (29, 28, 24) {real, imag} */,
  {32'h4245e309, 32'h4228c204} /* (29, 28, 23) {real, imag} */,
  {32'h4251e9e6, 32'h41fdc703} /* (29, 28, 22) {real, imag} */,
  {32'hc1dff779, 32'h423f9513} /* (29, 28, 21) {real, imag} */,
  {32'h4229abab, 32'hc1ab110c} /* (29, 28, 20) {real, imag} */,
  {32'h4143d7f8, 32'hc2692e54} /* (29, 28, 19) {real, imag} */,
  {32'h42b59938, 32'h4284232b} /* (29, 28, 18) {real, imag} */,
  {32'h401dbb22, 32'hc0fc2db6} /* (29, 28, 17) {real, imag} */,
  {32'h424ab333, 32'h00000000} /* (29, 28, 16) {real, imag} */,
  {32'h401dbb22, 32'h40fc2db6} /* (29, 28, 15) {real, imag} */,
  {32'h42b59938, 32'hc284232b} /* (29, 28, 14) {real, imag} */,
  {32'h4143d7f8, 32'h42692e54} /* (29, 28, 13) {real, imag} */,
  {32'h4229abab, 32'h41ab110c} /* (29, 28, 12) {real, imag} */,
  {32'hc1dff779, 32'hc23f9513} /* (29, 28, 11) {real, imag} */,
  {32'h4251e9e6, 32'hc1fdc703} /* (29, 28, 10) {real, imag} */,
  {32'h4245e309, 32'hc228c204} /* (29, 28, 9) {real, imag} */,
  {32'hc09a5af0, 32'hc23d77fc} /* (29, 28, 8) {real, imag} */,
  {32'hc2ce4658, 32'h428dde02} /* (29, 28, 7) {real, imag} */,
  {32'h423b1904, 32'h428315fb} /* (29, 28, 6) {real, imag} */,
  {32'hc34b8a56, 32'hc2d915de} /* (29, 28, 5) {real, imag} */,
  {32'h43593aca, 32'h4249ae6c} /* (29, 28, 4) {real, imag} */,
  {32'hc0acd4a8, 32'h43834130} /* (29, 28, 3) {real, imag} */,
  {32'hc48c409c, 32'hc39a1c8c} /* (29, 28, 2) {real, imag} */,
  {32'h44cae112, 32'h42c14650} /* (29, 28, 1) {real, imag} */,
  {32'h445479fb, 32'h00000000} /* (29, 28, 0) {real, imag} */,
  {32'h44d16735, 32'h426d2620} /* (29, 27, 31) {real, imag} */,
  {32'hc4a09dae, 32'h437358dc} /* (29, 27, 30) {real, imag} */,
  {32'hc2bb4225, 32'hc3028a7a} /* (29, 27, 29) {real, imag} */,
  {32'h435d8032, 32'hc13a681e} /* (29, 27, 28) {real, imag} */,
  {32'hc33a61e6, 32'h4302d3aa} /* (29, 27, 27) {real, imag} */,
  {32'h42944ae4, 32'hc280c477} /* (29, 27, 26) {real, imag} */,
  {32'hc2de821c, 32'hc3069df3} /* (29, 27, 25) {real, imag} */,
  {32'hc212993e, 32'h422e6f80} /* (29, 27, 24) {real, imag} */,
  {32'h4204f61e, 32'hc2649748} /* (29, 27, 23) {real, imag} */,
  {32'hc19735e0, 32'hc29e4387} /* (29, 27, 22) {real, imag} */,
  {32'h4284f248, 32'h4294a0fc} /* (29, 27, 21) {real, imag} */,
  {32'h412778f4, 32'h42a2c654} /* (29, 27, 20) {real, imag} */,
  {32'h4284908b, 32'h4211bc59} /* (29, 27, 19) {real, imag} */,
  {32'hc1a36d02, 32'h4189c72c} /* (29, 27, 18) {real, imag} */,
  {32'hc263dfdc, 32'h4003d220} /* (29, 27, 17) {real, imag} */,
  {32'hc211d460, 32'h00000000} /* (29, 27, 16) {real, imag} */,
  {32'hc263dfdc, 32'hc003d220} /* (29, 27, 15) {real, imag} */,
  {32'hc1a36d02, 32'hc189c72c} /* (29, 27, 14) {real, imag} */,
  {32'h4284908b, 32'hc211bc59} /* (29, 27, 13) {real, imag} */,
  {32'h412778f4, 32'hc2a2c654} /* (29, 27, 12) {real, imag} */,
  {32'h4284f248, 32'hc294a0fc} /* (29, 27, 11) {real, imag} */,
  {32'hc19735e0, 32'h429e4387} /* (29, 27, 10) {real, imag} */,
  {32'h4204f61e, 32'h42649748} /* (29, 27, 9) {real, imag} */,
  {32'hc212993e, 32'hc22e6f80} /* (29, 27, 8) {real, imag} */,
  {32'hc2de821c, 32'h43069df3} /* (29, 27, 7) {real, imag} */,
  {32'h42944ae4, 32'h4280c477} /* (29, 27, 6) {real, imag} */,
  {32'hc33a61e6, 32'hc302d3aa} /* (29, 27, 5) {real, imag} */,
  {32'h435d8032, 32'h413a681e} /* (29, 27, 4) {real, imag} */,
  {32'hc2bb4225, 32'h43028a7a} /* (29, 27, 3) {real, imag} */,
  {32'hc4a09dae, 32'hc37358dc} /* (29, 27, 2) {real, imag} */,
  {32'h44d16735, 32'hc26d2620} /* (29, 27, 1) {real, imag} */,
  {32'h4485efa3, 32'h00000000} /* (29, 27, 0) {real, imag} */,
  {32'h44d7a119, 32'hc1a3f9c0} /* (29, 26, 31) {real, imag} */,
  {32'hc494dd02, 32'h434da46c} /* (29, 26, 30) {real, imag} */,
  {32'hc29e90a2, 32'hc246d657} /* (29, 26, 29) {real, imag} */,
  {32'h42ecbf1e, 32'hc0618080} /* (29, 26, 28) {real, imag} */,
  {32'hc3341fac, 32'h41f79554} /* (29, 26, 27) {real, imag} */,
  {32'hc211a991, 32'h41a9cfb4} /* (29, 26, 26) {real, imag} */,
  {32'h421beb30, 32'hc20cc3ce} /* (29, 26, 25) {real, imag} */,
  {32'h410173bc, 32'h411f7d88} /* (29, 26, 24) {real, imag} */,
  {32'h4272556f, 32'hc1ebb39a} /* (29, 26, 23) {real, imag} */,
  {32'hc1657c1b, 32'h42038178} /* (29, 26, 22) {real, imag} */,
  {32'h42919fa4, 32'h41a86f6a} /* (29, 26, 21) {real, imag} */,
  {32'h42e3bc08, 32'hc13c74ca} /* (29, 26, 20) {real, imag} */,
  {32'hc1abeb60, 32'hc20fdb50} /* (29, 26, 19) {real, imag} */,
  {32'hc1f43e4c, 32'h41c8e4dc} /* (29, 26, 18) {real, imag} */,
  {32'h41077510, 32'h41f946a8} /* (29, 26, 17) {real, imag} */,
  {32'hc29d7199, 32'h00000000} /* (29, 26, 16) {real, imag} */,
  {32'h41077510, 32'hc1f946a8} /* (29, 26, 15) {real, imag} */,
  {32'hc1f43e4c, 32'hc1c8e4dc} /* (29, 26, 14) {real, imag} */,
  {32'hc1abeb60, 32'h420fdb50} /* (29, 26, 13) {real, imag} */,
  {32'h42e3bc08, 32'h413c74ca} /* (29, 26, 12) {real, imag} */,
  {32'h42919fa4, 32'hc1a86f6a} /* (29, 26, 11) {real, imag} */,
  {32'hc1657c1b, 32'hc2038178} /* (29, 26, 10) {real, imag} */,
  {32'h4272556f, 32'h41ebb39a} /* (29, 26, 9) {real, imag} */,
  {32'h410173bc, 32'hc11f7d88} /* (29, 26, 8) {real, imag} */,
  {32'h421beb30, 32'h420cc3ce} /* (29, 26, 7) {real, imag} */,
  {32'hc211a991, 32'hc1a9cfb4} /* (29, 26, 6) {real, imag} */,
  {32'hc3341fac, 32'hc1f79554} /* (29, 26, 5) {real, imag} */,
  {32'h42ecbf1e, 32'h40618080} /* (29, 26, 4) {real, imag} */,
  {32'hc29e90a2, 32'h4246d657} /* (29, 26, 3) {real, imag} */,
  {32'hc494dd02, 32'hc34da46c} /* (29, 26, 2) {real, imag} */,
  {32'h44d7a119, 32'h41a3f9c0} /* (29, 26, 1) {real, imag} */,
  {32'h4463d032, 32'h00000000} /* (29, 26, 0) {real, imag} */,
  {32'h44d39b92, 32'hc2bebe30} /* (29, 25, 31) {real, imag} */,
  {32'hc49907a6, 32'h438ee525} /* (29, 25, 30) {real, imag} */,
  {32'hc2b58dd4, 32'hc338a05a} /* (29, 25, 29) {real, imag} */,
  {32'h43217aa6, 32'h41a941c9} /* (29, 25, 28) {real, imag} */,
  {32'hc317a475, 32'hc1b42d72} /* (29, 25, 27) {real, imag} */,
  {32'h41d6dc76, 32'hc0e98078} /* (29, 25, 26) {real, imag} */,
  {32'hc1318340, 32'hc309a476} /* (29, 25, 25) {real, imag} */,
  {32'h4282b3e2, 32'h42895083} /* (29, 25, 24) {real, imag} */,
  {32'hc2864b86, 32'h4281ca2d} /* (29, 25, 23) {real, imag} */,
  {32'h429b7503, 32'hc1291d16} /* (29, 25, 22) {real, imag} */,
  {32'hc1849de0, 32'h41d92628} /* (29, 25, 21) {real, imag} */,
  {32'hc2335672, 32'h41bca24e} /* (29, 25, 20) {real, imag} */,
  {32'hc2478944, 32'hc2d120b3} /* (29, 25, 19) {real, imag} */,
  {32'hc151e9c0, 32'hc10e3590} /* (29, 25, 18) {real, imag} */,
  {32'h4205eae3, 32'hc25efb8c} /* (29, 25, 17) {real, imag} */,
  {32'h41281a2c, 32'h00000000} /* (29, 25, 16) {real, imag} */,
  {32'h4205eae3, 32'h425efb8c} /* (29, 25, 15) {real, imag} */,
  {32'hc151e9c0, 32'h410e3590} /* (29, 25, 14) {real, imag} */,
  {32'hc2478944, 32'h42d120b3} /* (29, 25, 13) {real, imag} */,
  {32'hc2335672, 32'hc1bca24e} /* (29, 25, 12) {real, imag} */,
  {32'hc1849de0, 32'hc1d92628} /* (29, 25, 11) {real, imag} */,
  {32'h429b7503, 32'h41291d16} /* (29, 25, 10) {real, imag} */,
  {32'hc2864b86, 32'hc281ca2d} /* (29, 25, 9) {real, imag} */,
  {32'h4282b3e2, 32'hc2895083} /* (29, 25, 8) {real, imag} */,
  {32'hc1318340, 32'h4309a476} /* (29, 25, 7) {real, imag} */,
  {32'h41d6dc76, 32'h40e98078} /* (29, 25, 6) {real, imag} */,
  {32'hc317a475, 32'h41b42d72} /* (29, 25, 5) {real, imag} */,
  {32'h43217aa6, 32'hc1a941c9} /* (29, 25, 4) {real, imag} */,
  {32'hc2b58dd4, 32'h4338a05a} /* (29, 25, 3) {real, imag} */,
  {32'hc49907a6, 32'hc38ee525} /* (29, 25, 2) {real, imag} */,
  {32'h44d39b92, 32'h42bebe30} /* (29, 25, 1) {real, imag} */,
  {32'h44671a75, 32'h00000000} /* (29, 25, 0) {real, imag} */,
  {32'h44ca382e, 32'h41e47380} /* (29, 24, 31) {real, imag} */,
  {32'hc4a52f32, 32'h43976100} /* (29, 24, 30) {real, imag} */,
  {32'hc22cc8f3, 32'h40d58a56} /* (29, 24, 29) {real, imag} */,
  {32'h438a3a4a, 32'hc19d89b8} /* (29, 24, 28) {real, imag} */,
  {32'hc2460d54, 32'h42809ee2} /* (29, 24, 27) {real, imag} */,
  {32'hc1da5384, 32'hbf89eec0} /* (29, 24, 26) {real, imag} */,
  {32'hc323501a, 32'hc2dc37e4} /* (29, 24, 25) {real, imag} */,
  {32'hc28a0fa1, 32'h424b3c9e} /* (29, 24, 24) {real, imag} */,
  {32'hc1bd8c2f, 32'hc2313d7a} /* (29, 24, 23) {real, imag} */,
  {32'hbfba2580, 32'hc3197aac} /* (29, 24, 22) {real, imag} */,
  {32'hc2034c74, 32'h427fcf15} /* (29, 24, 21) {real, imag} */,
  {32'hc1abdd9e, 32'h41eae93e} /* (29, 24, 20) {real, imag} */,
  {32'h41a92bd9, 32'h42303ca8} /* (29, 24, 19) {real, imag} */,
  {32'h40a76e20, 32'h42073bd0} /* (29, 24, 18) {real, imag} */,
  {32'h4283424f, 32'hc281e2a0} /* (29, 24, 17) {real, imag} */,
  {32'hc18ff57a, 32'h00000000} /* (29, 24, 16) {real, imag} */,
  {32'h4283424f, 32'h4281e2a0} /* (29, 24, 15) {real, imag} */,
  {32'h40a76e20, 32'hc2073bd0} /* (29, 24, 14) {real, imag} */,
  {32'h41a92bd9, 32'hc2303ca8} /* (29, 24, 13) {real, imag} */,
  {32'hc1abdd9e, 32'hc1eae93e} /* (29, 24, 12) {real, imag} */,
  {32'hc2034c74, 32'hc27fcf15} /* (29, 24, 11) {real, imag} */,
  {32'hbfba2580, 32'h43197aac} /* (29, 24, 10) {real, imag} */,
  {32'hc1bd8c2f, 32'h42313d7a} /* (29, 24, 9) {real, imag} */,
  {32'hc28a0fa1, 32'hc24b3c9e} /* (29, 24, 8) {real, imag} */,
  {32'hc323501a, 32'h42dc37e4} /* (29, 24, 7) {real, imag} */,
  {32'hc1da5384, 32'h3f89eec0} /* (29, 24, 6) {real, imag} */,
  {32'hc2460d54, 32'hc2809ee2} /* (29, 24, 5) {real, imag} */,
  {32'h438a3a4a, 32'h419d89b8} /* (29, 24, 4) {real, imag} */,
  {32'hc22cc8f3, 32'hc0d58a56} /* (29, 24, 3) {real, imag} */,
  {32'hc4a52f32, 32'hc3976100} /* (29, 24, 2) {real, imag} */,
  {32'h44ca382e, 32'hc1e47380} /* (29, 24, 1) {real, imag} */,
  {32'h448632e0, 32'h00000000} /* (29, 24, 0) {real, imag} */,
  {32'h44a2ce2a, 32'h42d7c63c} /* (29, 23, 31) {real, imag} */,
  {32'hc476a35e, 32'h4375ead2} /* (29, 23, 30) {real, imag} */,
  {32'hc196e636, 32'h4290ad77} /* (29, 23, 29) {real, imag} */,
  {32'h42ee87c6, 32'hc322ea03} /* (29, 23, 28) {real, imag} */,
  {32'hc2a16afa, 32'h430b71c6} /* (29, 23, 27) {real, imag} */,
  {32'h425b9f75, 32'hc2576fa5} /* (29, 23, 26) {real, imag} */,
  {32'hc302c16e, 32'hc2f0c9f2} /* (29, 23, 25) {real, imag} */,
  {32'hc163c4a6, 32'h413fe8a2} /* (29, 23, 24) {real, imag} */,
  {32'hc19a270c, 32'h420fd621} /* (29, 23, 23) {real, imag} */,
  {32'h4264aac4, 32'h4182b148} /* (29, 23, 22) {real, imag} */,
  {32'h3f34f800, 32'hc2c0c5a9} /* (29, 23, 21) {real, imag} */,
  {32'hc19aea8a, 32'h41a1dacc} /* (29, 23, 20) {real, imag} */,
  {32'hc1516b0e, 32'hc09dc88e} /* (29, 23, 19) {real, imag} */,
  {32'hc2ecb644, 32'h41d9e2c0} /* (29, 23, 18) {real, imag} */,
  {32'h41acf5ca, 32'hc17412dc} /* (29, 23, 17) {real, imag} */,
  {32'hc2882122, 32'h00000000} /* (29, 23, 16) {real, imag} */,
  {32'h41acf5ca, 32'h417412dc} /* (29, 23, 15) {real, imag} */,
  {32'hc2ecb644, 32'hc1d9e2c0} /* (29, 23, 14) {real, imag} */,
  {32'hc1516b0e, 32'h409dc88e} /* (29, 23, 13) {real, imag} */,
  {32'hc19aea8a, 32'hc1a1dacc} /* (29, 23, 12) {real, imag} */,
  {32'h3f34f800, 32'h42c0c5a9} /* (29, 23, 11) {real, imag} */,
  {32'h4264aac4, 32'hc182b148} /* (29, 23, 10) {real, imag} */,
  {32'hc19a270c, 32'hc20fd621} /* (29, 23, 9) {real, imag} */,
  {32'hc163c4a6, 32'hc13fe8a2} /* (29, 23, 8) {real, imag} */,
  {32'hc302c16e, 32'h42f0c9f2} /* (29, 23, 7) {real, imag} */,
  {32'h425b9f75, 32'h42576fa5} /* (29, 23, 6) {real, imag} */,
  {32'hc2a16afa, 32'hc30b71c6} /* (29, 23, 5) {real, imag} */,
  {32'h42ee87c6, 32'h4322ea03} /* (29, 23, 4) {real, imag} */,
  {32'hc196e636, 32'hc290ad77} /* (29, 23, 3) {real, imag} */,
  {32'hc476a35e, 32'hc375ead2} /* (29, 23, 2) {real, imag} */,
  {32'h44a2ce2a, 32'hc2d7c63c} /* (29, 23, 1) {real, imag} */,
  {32'h445a93b0, 32'h00000000} /* (29, 23, 0) {real, imag} */,
  {32'h44574720, 32'h42328392} /* (29, 22, 31) {real, imag} */,
  {32'hc408deb6, 32'h43a8a094} /* (29, 22, 30) {real, imag} */,
  {32'h3e2b3e00, 32'h42ec719f} /* (29, 22, 29) {real, imag} */,
  {32'h4300d624, 32'hc22fad4c} /* (29, 22, 28) {real, imag} */,
  {32'hc2d807f5, 32'h4260a7a9} /* (29, 22, 27) {real, imag} */,
  {32'hc0399d30, 32'h42c300b4} /* (29, 22, 26) {real, imag} */,
  {32'h40251a20, 32'hc009e3a8} /* (29, 22, 25) {real, imag} */,
  {32'hc2cd5bc8, 32'h417662d8} /* (29, 22, 24) {real, imag} */,
  {32'h4071a2d8, 32'h426b4bd1} /* (29, 22, 23) {real, imag} */,
  {32'hc14ef357, 32'hc24b40e8} /* (29, 22, 22) {real, imag} */,
  {32'hc251fb5f, 32'hc1e07448} /* (29, 22, 21) {real, imag} */,
  {32'h3febbf80, 32'hc2e11e6a} /* (29, 22, 20) {real, imag} */,
  {32'hc286e720, 32'hc28d90ce} /* (29, 22, 19) {real, imag} */,
  {32'hc1a48168, 32'h42c72fad} /* (29, 22, 18) {real, imag} */,
  {32'h4017db72, 32'hc2367810} /* (29, 22, 17) {real, imag} */,
  {32'hc24700c5, 32'h00000000} /* (29, 22, 16) {real, imag} */,
  {32'h4017db72, 32'h42367810} /* (29, 22, 15) {real, imag} */,
  {32'hc1a48168, 32'hc2c72fad} /* (29, 22, 14) {real, imag} */,
  {32'hc286e720, 32'h428d90ce} /* (29, 22, 13) {real, imag} */,
  {32'h3febbf80, 32'h42e11e6a} /* (29, 22, 12) {real, imag} */,
  {32'hc251fb5f, 32'h41e07448} /* (29, 22, 11) {real, imag} */,
  {32'hc14ef357, 32'h424b40e8} /* (29, 22, 10) {real, imag} */,
  {32'h4071a2d8, 32'hc26b4bd1} /* (29, 22, 9) {real, imag} */,
  {32'hc2cd5bc8, 32'hc17662d8} /* (29, 22, 8) {real, imag} */,
  {32'h40251a20, 32'h4009e3a8} /* (29, 22, 7) {real, imag} */,
  {32'hc0399d30, 32'hc2c300b4} /* (29, 22, 6) {real, imag} */,
  {32'hc2d807f5, 32'hc260a7a9} /* (29, 22, 5) {real, imag} */,
  {32'h4300d624, 32'h422fad4c} /* (29, 22, 4) {real, imag} */,
  {32'h3e2b3e00, 32'hc2ec719f} /* (29, 22, 3) {real, imag} */,
  {32'hc408deb6, 32'hc3a8a094} /* (29, 22, 2) {real, imag} */,
  {32'h44574720, 32'hc2328392} /* (29, 22, 1) {real, imag} */,
  {32'h443eaf6a, 32'h00000000} /* (29, 22, 0) {real, imag} */,
  {32'h41edcce0, 32'h431c67a9} /* (29, 21, 31) {real, imag} */,
  {32'hc320d0e2, 32'hc03c20c0} /* (29, 21, 30) {real, imag} */,
  {32'h436c8412, 32'hc1d746be} /* (29, 21, 29) {real, imag} */,
  {32'hc18f1908, 32'h42193122} /* (29, 21, 28) {real, imag} */,
  {32'hc2875b40, 32'hc2930abc} /* (29, 21, 27) {real, imag} */,
  {32'hc27e70d6, 32'h42904ef3} /* (29, 21, 26) {real, imag} */,
  {32'hc2939a10, 32'hc1fc14c2} /* (29, 21, 25) {real, imag} */,
  {32'h416517e8, 32'h41f0fef2} /* (29, 21, 24) {real, imag} */,
  {32'h41e11733, 32'hc2372d3e} /* (29, 21, 23) {real, imag} */,
  {32'hc1659659, 32'hbf28bfa0} /* (29, 21, 22) {real, imag} */,
  {32'hc23c7b58, 32'h42cb9c54} /* (29, 21, 21) {real, imag} */,
  {32'h41a3a28a, 32'hc18dee18} /* (29, 21, 20) {real, imag} */,
  {32'h42051ad1, 32'hc2a3b696} /* (29, 21, 19) {real, imag} */,
  {32'h41bae354, 32'h41155e1e} /* (29, 21, 18) {real, imag} */,
  {32'hc2382f88, 32'h42516944} /* (29, 21, 17) {real, imag} */,
  {32'h41fd2d2c, 32'h00000000} /* (29, 21, 16) {real, imag} */,
  {32'hc2382f88, 32'hc2516944} /* (29, 21, 15) {real, imag} */,
  {32'h41bae354, 32'hc1155e1e} /* (29, 21, 14) {real, imag} */,
  {32'h42051ad1, 32'h42a3b696} /* (29, 21, 13) {real, imag} */,
  {32'h41a3a28a, 32'h418dee18} /* (29, 21, 12) {real, imag} */,
  {32'hc23c7b58, 32'hc2cb9c54} /* (29, 21, 11) {real, imag} */,
  {32'hc1659659, 32'h3f28bfa0} /* (29, 21, 10) {real, imag} */,
  {32'h41e11733, 32'h42372d3e} /* (29, 21, 9) {real, imag} */,
  {32'h416517e8, 32'hc1f0fef2} /* (29, 21, 8) {real, imag} */,
  {32'hc2939a10, 32'h41fc14c2} /* (29, 21, 7) {real, imag} */,
  {32'hc27e70d6, 32'hc2904ef3} /* (29, 21, 6) {real, imag} */,
  {32'hc2875b40, 32'h42930abc} /* (29, 21, 5) {real, imag} */,
  {32'hc18f1908, 32'hc2193122} /* (29, 21, 4) {real, imag} */,
  {32'h436c8412, 32'h41d746be} /* (29, 21, 3) {real, imag} */,
  {32'hc320d0e2, 32'h403c20c0} /* (29, 21, 2) {real, imag} */,
  {32'h41edcce0, 32'hc31c67a9} /* (29, 21, 1) {real, imag} */,
  {32'h4202dc38, 32'h00000000} /* (29, 21, 0) {real, imag} */,
  {32'hc4921729, 32'h430c3b3a} /* (29, 20, 31) {real, imag} */,
  {32'h43ec5354, 32'hc3522cda} /* (29, 20, 30) {real, imag} */,
  {32'h432cda50, 32'hc2ba58e0} /* (29, 20, 29) {real, imag} */,
  {32'hc21d5f46, 32'hc1d47822} /* (29, 20, 28) {real, imag} */,
  {32'h43266592, 32'hc265d79c} /* (29, 20, 27) {real, imag} */,
  {32'h407e5000, 32'hc21a5ade} /* (29, 20, 26) {real, imag} */,
  {32'h421618da, 32'hc28f6420} /* (29, 20, 25) {real, imag} */,
  {32'h42133064, 32'hbf5c2700} /* (29, 20, 24) {real, imag} */,
  {32'h422b2bfb, 32'h429021bc} /* (29, 20, 23) {real, imag} */,
  {32'hc19a39c0, 32'h42e046b3} /* (29, 20, 22) {real, imag} */,
  {32'hc2029965, 32'h41ae269e} /* (29, 20, 21) {real, imag} */,
  {32'hbe09fe00, 32'hc1c88e24} /* (29, 20, 20) {real, imag} */,
  {32'h419bbf91, 32'h4167b07c} /* (29, 20, 19) {real, imag} */,
  {32'h424dbbf5, 32'hc2765d52} /* (29, 20, 18) {real, imag} */,
  {32'h41c686da, 32'hc1d1a30d} /* (29, 20, 17) {real, imag} */,
  {32'h41cd30f2, 32'h00000000} /* (29, 20, 16) {real, imag} */,
  {32'h41c686da, 32'h41d1a30d} /* (29, 20, 15) {real, imag} */,
  {32'h424dbbf5, 32'h42765d52} /* (29, 20, 14) {real, imag} */,
  {32'h419bbf91, 32'hc167b07c} /* (29, 20, 13) {real, imag} */,
  {32'hbe09fe00, 32'h41c88e24} /* (29, 20, 12) {real, imag} */,
  {32'hc2029965, 32'hc1ae269e} /* (29, 20, 11) {real, imag} */,
  {32'hc19a39c0, 32'hc2e046b3} /* (29, 20, 10) {real, imag} */,
  {32'h422b2bfb, 32'hc29021bc} /* (29, 20, 9) {real, imag} */,
  {32'h42133064, 32'h3f5c2700} /* (29, 20, 8) {real, imag} */,
  {32'h421618da, 32'h428f6420} /* (29, 20, 7) {real, imag} */,
  {32'h407e5000, 32'h421a5ade} /* (29, 20, 6) {real, imag} */,
  {32'h43266592, 32'h4265d79c} /* (29, 20, 5) {real, imag} */,
  {32'hc21d5f46, 32'h41d47822} /* (29, 20, 4) {real, imag} */,
  {32'h432cda50, 32'h42ba58e0} /* (29, 20, 3) {real, imag} */,
  {32'h43ec5354, 32'h43522cda} /* (29, 20, 2) {real, imag} */,
  {32'hc4921729, 32'hc30c3b3a} /* (29, 20, 1) {real, imag} */,
  {32'hc449d366, 32'h00000000} /* (29, 20, 0) {real, imag} */,
  {32'hc4d9eb0c, 32'h431d5264} /* (29, 19, 31) {real, imag} */,
  {32'h442a07c0, 32'hc3814b15} /* (29, 19, 30) {real, imag} */,
  {32'h421e1a54, 32'h42f68766} /* (29, 19, 29) {real, imag} */,
  {32'hc36320e5, 32'h42e54c10} /* (29, 19, 28) {real, imag} */,
  {32'h4356da7e, 32'hc30d4d4c} /* (29, 19, 27) {real, imag} */,
  {32'h421ca7ac, 32'hc280b600} /* (29, 19, 26) {real, imag} */,
  {32'hc263fb96, 32'h41f9396e} /* (29, 19, 25) {real, imag} */,
  {32'h42712cc2, 32'hc16f708c} /* (29, 19, 24) {real, imag} */,
  {32'hc2329eb0, 32'hc31749e8} /* (29, 19, 23) {real, imag} */,
  {32'h401a22b8, 32'h42938346} /* (29, 19, 22) {real, imag} */,
  {32'h430f562c, 32'h421a3a8c} /* (29, 19, 21) {real, imag} */,
  {32'h41e9e9e9, 32'h429037fa} /* (29, 19, 20) {real, imag} */,
  {32'hc2531efa, 32'h425d4500} /* (29, 19, 19) {real, imag} */,
  {32'h419cc444, 32'h42b598f3} /* (29, 19, 18) {real, imag} */,
  {32'h42981289, 32'h40b46cf6} /* (29, 19, 17) {real, imag} */,
  {32'h41c193be, 32'h00000000} /* (29, 19, 16) {real, imag} */,
  {32'h42981289, 32'hc0b46cf6} /* (29, 19, 15) {real, imag} */,
  {32'h419cc444, 32'hc2b598f3} /* (29, 19, 14) {real, imag} */,
  {32'hc2531efa, 32'hc25d4500} /* (29, 19, 13) {real, imag} */,
  {32'h41e9e9e9, 32'hc29037fa} /* (29, 19, 12) {real, imag} */,
  {32'h430f562c, 32'hc21a3a8c} /* (29, 19, 11) {real, imag} */,
  {32'h401a22b8, 32'hc2938346} /* (29, 19, 10) {real, imag} */,
  {32'hc2329eb0, 32'h431749e8} /* (29, 19, 9) {real, imag} */,
  {32'h42712cc2, 32'h416f708c} /* (29, 19, 8) {real, imag} */,
  {32'hc263fb96, 32'hc1f9396e} /* (29, 19, 7) {real, imag} */,
  {32'h421ca7ac, 32'h4280b600} /* (29, 19, 6) {real, imag} */,
  {32'h4356da7e, 32'h430d4d4c} /* (29, 19, 5) {real, imag} */,
  {32'hc36320e5, 32'hc2e54c10} /* (29, 19, 4) {real, imag} */,
  {32'h421e1a54, 32'hc2f68766} /* (29, 19, 3) {real, imag} */,
  {32'h442a07c0, 32'h43814b15} /* (29, 19, 2) {real, imag} */,
  {32'hc4d9eb0c, 32'hc31d5264} /* (29, 19, 1) {real, imag} */,
  {32'hc48aba4b, 32'h00000000} /* (29, 19, 0) {real, imag} */,
  {32'hc4ff1691, 32'h43698cbc} /* (29, 18, 31) {real, imag} */,
  {32'h44524b60, 32'hc35c0e04} /* (29, 18, 30) {real, imag} */,
  {32'hc2cfa414, 32'hc1b21764} /* (29, 18, 29) {real, imag} */,
  {32'hc3276999, 32'h42461ce6} /* (29, 18, 28) {real, imag} */,
  {32'h438148bd, 32'hc333965d} /* (29, 18, 27) {real, imag} */,
  {32'hc2ae142e, 32'h41c94320} /* (29, 18, 26) {real, imag} */,
  {32'hc2fac06a, 32'h42baf9b0} /* (29, 18, 25) {real, imag} */,
  {32'h4088b200, 32'hc2620d0a} /* (29, 18, 24) {real, imag} */,
  {32'h427fdc7c, 32'h423cb5b6} /* (29, 18, 23) {real, imag} */,
  {32'hc2ba65b9, 32'hc20e7a7e} /* (29, 18, 22) {real, imag} */,
  {32'hc24762b6, 32'h3fcf8240} /* (29, 18, 21) {real, imag} */,
  {32'h42357502, 32'hc284d870} /* (29, 18, 20) {real, imag} */,
  {32'hc0c1e8d0, 32'h423455e2} /* (29, 18, 19) {real, imag} */,
  {32'h41b7deb6, 32'hc1d5837d} /* (29, 18, 18) {real, imag} */,
  {32'hc25a8148, 32'h41d9ca2c} /* (29, 18, 17) {real, imag} */,
  {32'h42850449, 32'h00000000} /* (29, 18, 16) {real, imag} */,
  {32'hc25a8148, 32'hc1d9ca2c} /* (29, 18, 15) {real, imag} */,
  {32'h41b7deb6, 32'h41d5837d} /* (29, 18, 14) {real, imag} */,
  {32'hc0c1e8d0, 32'hc23455e2} /* (29, 18, 13) {real, imag} */,
  {32'h42357502, 32'h4284d870} /* (29, 18, 12) {real, imag} */,
  {32'hc24762b6, 32'hbfcf8240} /* (29, 18, 11) {real, imag} */,
  {32'hc2ba65b9, 32'h420e7a7e} /* (29, 18, 10) {real, imag} */,
  {32'h427fdc7c, 32'hc23cb5b6} /* (29, 18, 9) {real, imag} */,
  {32'h4088b200, 32'h42620d0a} /* (29, 18, 8) {real, imag} */,
  {32'hc2fac06a, 32'hc2baf9b0} /* (29, 18, 7) {real, imag} */,
  {32'hc2ae142e, 32'hc1c94320} /* (29, 18, 6) {real, imag} */,
  {32'h438148bd, 32'h4333965d} /* (29, 18, 5) {real, imag} */,
  {32'hc3276999, 32'hc2461ce6} /* (29, 18, 4) {real, imag} */,
  {32'hc2cfa414, 32'h41b21764} /* (29, 18, 3) {real, imag} */,
  {32'h44524b60, 32'h435c0e04} /* (29, 18, 2) {real, imag} */,
  {32'hc4ff1691, 32'hc3698cbc} /* (29, 18, 1) {real, imag} */,
  {32'hc4bf409e, 32'h00000000} /* (29, 18, 0) {real, imag} */,
  {32'hc503f884, 32'h43b51874} /* (29, 17, 31) {real, imag} */,
  {32'h447d692d, 32'hc344ec4e} /* (29, 17, 30) {real, imag} */,
  {32'hc2aedc81, 32'h42bbf7a3} /* (29, 17, 29) {real, imag} */,
  {32'h4191df28, 32'h42d85064} /* (29, 17, 28) {real, imag} */,
  {32'h4319f445, 32'hc32464aa} /* (29, 17, 27) {real, imag} */,
  {32'h41e3fe6c, 32'h3f81e670} /* (29, 17, 26) {real, imag} */,
  {32'h4281a2ae, 32'h429ae334} /* (29, 17, 25) {real, imag} */,
  {32'h41a97602, 32'h423595f7} /* (29, 17, 24) {real, imag} */,
  {32'h42350ed4, 32'hc135d736} /* (29, 17, 23) {real, imag} */,
  {32'h4181ed95, 32'h400f8558} /* (29, 17, 22) {real, imag} */,
  {32'h4221c177, 32'hc2b81252} /* (29, 17, 21) {real, imag} */,
  {32'hc20b99e2, 32'h4293ddb6} /* (29, 17, 20) {real, imag} */,
  {32'h42d8dca8, 32'hc309088f} /* (29, 17, 19) {real, imag} */,
  {32'hc1cd4e51, 32'hc148631c} /* (29, 17, 18) {real, imag} */,
  {32'hc21b577e, 32'hc22bbbfc} /* (29, 17, 17) {real, imag} */,
  {32'hc29b1c01, 32'h00000000} /* (29, 17, 16) {real, imag} */,
  {32'hc21b577e, 32'h422bbbfc} /* (29, 17, 15) {real, imag} */,
  {32'hc1cd4e51, 32'h4148631c} /* (29, 17, 14) {real, imag} */,
  {32'h42d8dca8, 32'h4309088f} /* (29, 17, 13) {real, imag} */,
  {32'hc20b99e2, 32'hc293ddb6} /* (29, 17, 12) {real, imag} */,
  {32'h4221c177, 32'h42b81252} /* (29, 17, 11) {real, imag} */,
  {32'h4181ed95, 32'hc00f8558} /* (29, 17, 10) {real, imag} */,
  {32'h42350ed4, 32'h4135d736} /* (29, 17, 9) {real, imag} */,
  {32'h41a97602, 32'hc23595f7} /* (29, 17, 8) {real, imag} */,
  {32'h4281a2ae, 32'hc29ae334} /* (29, 17, 7) {real, imag} */,
  {32'h41e3fe6c, 32'hbf81e670} /* (29, 17, 6) {real, imag} */,
  {32'h4319f445, 32'h432464aa} /* (29, 17, 5) {real, imag} */,
  {32'h4191df28, 32'hc2d85064} /* (29, 17, 4) {real, imag} */,
  {32'hc2aedc81, 32'hc2bbf7a3} /* (29, 17, 3) {real, imag} */,
  {32'h447d692d, 32'h4344ec4e} /* (29, 17, 2) {real, imag} */,
  {32'hc503f884, 32'hc3b51874} /* (29, 17, 1) {real, imag} */,
  {32'hc4d71924, 32'h00000000} /* (29, 17, 0) {real, imag} */,
  {32'hc5041544, 32'h434878c0} /* (29, 16, 31) {real, imag} */,
  {32'h4480bc8d, 32'hc3548854} /* (29, 16, 30) {real, imag} */,
  {32'hc25e1ca2, 32'h4225569a} /* (29, 16, 29) {real, imag} */,
  {32'hc2854d6e, 32'h423369f0} /* (29, 16, 28) {real, imag} */,
  {32'h4304350b, 32'hc299d78c} /* (29, 16, 27) {real, imag} */,
  {32'h42552700, 32'hc2e97066} /* (29, 16, 26) {real, imag} */,
  {32'hbfceb830, 32'h42669506} /* (29, 16, 25) {real, imag} */,
  {32'hc1209f8b, 32'hc21de6b8} /* (29, 16, 24) {real, imag} */,
  {32'hbf1413e0, 32'h42026fe8} /* (29, 16, 23) {real, imag} */,
  {32'h430b3037, 32'hc1b84003} /* (29, 16, 22) {real, imag} */,
  {32'h41d60336, 32'hc2ff448b} /* (29, 16, 21) {real, imag} */,
  {32'hc2af3dfc, 32'hc2b7203a} /* (29, 16, 20) {real, imag} */,
  {32'h417a2fa2, 32'hc27c12fa} /* (29, 16, 19) {real, imag} */,
  {32'h41b792a0, 32'hc1b4f8db} /* (29, 16, 18) {real, imag} */,
  {32'h4238eff8, 32'h429c1f42} /* (29, 16, 17) {real, imag} */,
  {32'h40a6d684, 32'h00000000} /* (29, 16, 16) {real, imag} */,
  {32'h4238eff8, 32'hc29c1f42} /* (29, 16, 15) {real, imag} */,
  {32'h41b792a0, 32'h41b4f8db} /* (29, 16, 14) {real, imag} */,
  {32'h417a2fa2, 32'h427c12fa} /* (29, 16, 13) {real, imag} */,
  {32'hc2af3dfc, 32'h42b7203a} /* (29, 16, 12) {real, imag} */,
  {32'h41d60336, 32'h42ff448b} /* (29, 16, 11) {real, imag} */,
  {32'h430b3037, 32'h41b84003} /* (29, 16, 10) {real, imag} */,
  {32'hbf1413e0, 32'hc2026fe8} /* (29, 16, 9) {real, imag} */,
  {32'hc1209f8b, 32'h421de6b8} /* (29, 16, 8) {real, imag} */,
  {32'hbfceb830, 32'hc2669506} /* (29, 16, 7) {real, imag} */,
  {32'h42552700, 32'h42e97066} /* (29, 16, 6) {real, imag} */,
  {32'h4304350b, 32'h4299d78c} /* (29, 16, 5) {real, imag} */,
  {32'hc2854d6e, 32'hc23369f0} /* (29, 16, 4) {real, imag} */,
  {32'hc25e1ca2, 32'hc225569a} /* (29, 16, 3) {real, imag} */,
  {32'h4480bc8d, 32'h43548854} /* (29, 16, 2) {real, imag} */,
  {32'hc5041544, 32'hc34878c0} /* (29, 16, 1) {real, imag} */,
  {32'hc4d97e25, 32'h00000000} /* (29, 16, 0) {real, imag} */,
  {32'hc4fd72dd, 32'h41c4a3c8} /* (29, 15, 31) {real, imag} */,
  {32'h44897c78, 32'hc3680632} /* (29, 15, 30) {real, imag} */,
  {32'h418973e8, 32'h4349abaa} /* (29, 15, 29) {real, imag} */,
  {32'hc35b1381, 32'h40f3ace0} /* (29, 15, 28) {real, imag} */,
  {32'h428315f8, 32'h41db98a0} /* (29, 15, 27) {real, imag} */,
  {32'h4282dfff, 32'hc22ad1d0} /* (29, 15, 26) {real, imag} */,
  {32'h427488a8, 32'h4193783e} /* (29, 15, 25) {real, imag} */,
  {32'h42d5763a, 32'hc22405ed} /* (29, 15, 24) {real, imag} */,
  {32'hc2a2ac9c, 32'h41ff1985} /* (29, 15, 23) {real, imag} */,
  {32'hc1131ba2, 32'hc27813ce} /* (29, 15, 22) {real, imag} */,
  {32'h430740d6, 32'hc138b7a4} /* (29, 15, 21) {real, imag} */,
  {32'h41630481, 32'h418ee6d0} /* (29, 15, 20) {real, imag} */,
  {32'hc28780d0, 32'h4247521c} /* (29, 15, 19) {real, imag} */,
  {32'hc171944a, 32'hc27439ef} /* (29, 15, 18) {real, imag} */,
  {32'hc2598598, 32'hc1fd4664} /* (29, 15, 17) {real, imag} */,
  {32'h42d24b2b, 32'h00000000} /* (29, 15, 16) {real, imag} */,
  {32'hc2598598, 32'h41fd4664} /* (29, 15, 15) {real, imag} */,
  {32'hc171944a, 32'h427439ef} /* (29, 15, 14) {real, imag} */,
  {32'hc28780d0, 32'hc247521c} /* (29, 15, 13) {real, imag} */,
  {32'h41630481, 32'hc18ee6d0} /* (29, 15, 12) {real, imag} */,
  {32'h430740d6, 32'h4138b7a4} /* (29, 15, 11) {real, imag} */,
  {32'hc1131ba2, 32'h427813ce} /* (29, 15, 10) {real, imag} */,
  {32'hc2a2ac9c, 32'hc1ff1985} /* (29, 15, 9) {real, imag} */,
  {32'h42d5763a, 32'h422405ed} /* (29, 15, 8) {real, imag} */,
  {32'h427488a8, 32'hc193783e} /* (29, 15, 7) {real, imag} */,
  {32'h4282dfff, 32'h422ad1d0} /* (29, 15, 6) {real, imag} */,
  {32'h428315f8, 32'hc1db98a0} /* (29, 15, 5) {real, imag} */,
  {32'hc35b1381, 32'hc0f3ace0} /* (29, 15, 4) {real, imag} */,
  {32'h418973e8, 32'hc349abaa} /* (29, 15, 3) {real, imag} */,
  {32'h44897c78, 32'h43680632} /* (29, 15, 2) {real, imag} */,
  {32'hc4fd72dd, 32'hc1c4a3c8} /* (29, 15, 1) {real, imag} */,
  {32'hc4be78c8, 32'h00000000} /* (29, 15, 0) {real, imag} */,
  {32'hc4f2a10b, 32'h43129de8} /* (29, 14, 31) {real, imag} */,
  {32'h44821706, 32'hc384f118} /* (29, 14, 30) {real, imag} */,
  {32'hc28a6f42, 32'h42bdafef} /* (29, 14, 29) {real, imag} */,
  {32'hc354c12d, 32'h42fa9a0d} /* (29, 14, 28) {real, imag} */,
  {32'h43568b3f, 32'h41f02478} /* (29, 14, 27) {real, imag} */,
  {32'h4324dd13, 32'hc1b43188} /* (29, 14, 26) {real, imag} */,
  {32'hc2614b94, 32'h42656fff} /* (29, 14, 25) {real, imag} */,
  {32'h42a4dd22, 32'hc29649bd} /* (29, 14, 24) {real, imag} */,
  {32'h42869aea, 32'h412624ec} /* (29, 14, 23) {real, imag} */,
  {32'hc24f489e, 32'h42f094b3} /* (29, 14, 22) {real, imag} */,
  {32'hc2154c8e, 32'hc2ba3261} /* (29, 14, 21) {real, imag} */,
  {32'hc2b4cead, 32'h42227b34} /* (29, 14, 20) {real, imag} */,
  {32'hc2c0f595, 32'h417238b6} /* (29, 14, 19) {real, imag} */,
  {32'hc07bdf34, 32'h40cb3fac} /* (29, 14, 18) {real, imag} */,
  {32'hc197ea10, 32'hc2baaafb} /* (29, 14, 17) {real, imag} */,
  {32'h428bd94b, 32'h00000000} /* (29, 14, 16) {real, imag} */,
  {32'hc197ea10, 32'h42baaafb} /* (29, 14, 15) {real, imag} */,
  {32'hc07bdf34, 32'hc0cb3fac} /* (29, 14, 14) {real, imag} */,
  {32'hc2c0f595, 32'hc17238b6} /* (29, 14, 13) {real, imag} */,
  {32'hc2b4cead, 32'hc2227b34} /* (29, 14, 12) {real, imag} */,
  {32'hc2154c8e, 32'h42ba3261} /* (29, 14, 11) {real, imag} */,
  {32'hc24f489e, 32'hc2f094b3} /* (29, 14, 10) {real, imag} */,
  {32'h42869aea, 32'hc12624ec} /* (29, 14, 9) {real, imag} */,
  {32'h42a4dd22, 32'h429649bd} /* (29, 14, 8) {real, imag} */,
  {32'hc2614b94, 32'hc2656fff} /* (29, 14, 7) {real, imag} */,
  {32'h4324dd13, 32'h41b43188} /* (29, 14, 6) {real, imag} */,
  {32'h43568b3f, 32'hc1f02478} /* (29, 14, 5) {real, imag} */,
  {32'hc354c12d, 32'hc2fa9a0d} /* (29, 14, 4) {real, imag} */,
  {32'hc28a6f42, 32'hc2bdafef} /* (29, 14, 3) {real, imag} */,
  {32'h44821706, 32'h4384f118} /* (29, 14, 2) {real, imag} */,
  {32'hc4f2a10b, 32'hc3129de8} /* (29, 14, 1) {real, imag} */,
  {32'hc4c4df0e, 32'h00000000} /* (29, 14, 0) {real, imag} */,
  {32'hc4e1bee2, 32'h432a7014} /* (29, 13, 31) {real, imag} */,
  {32'h4474df0c, 32'hc31d230a} /* (29, 13, 30) {real, imag} */,
  {32'hc242621c, 32'hc20eb58f} /* (29, 13, 29) {real, imag} */,
  {32'hc3531b27, 32'h42ee22ec} /* (29, 13, 28) {real, imag} */,
  {32'h438cd8e1, 32'hc31775b4} /* (29, 13, 27) {real, imag} */,
  {32'h42e60748, 32'h42e94ffe} /* (29, 13, 26) {real, imag} */,
  {32'hc0b910cc, 32'h41b1e822} /* (29, 13, 25) {real, imag} */,
  {32'hc127f05a, 32'hc2d097a4} /* (29, 13, 24) {real, imag} */,
  {32'hc2d76482, 32'h42c24a86} /* (29, 13, 23) {real, imag} */,
  {32'h42768b20, 32'h422573d9} /* (29, 13, 22) {real, imag} */,
  {32'h423a95e7, 32'h427d31bc} /* (29, 13, 21) {real, imag} */,
  {32'hc1946cc1, 32'hc14dfb98} /* (29, 13, 20) {real, imag} */,
  {32'hc26c3b6e, 32'hc244a7a4} /* (29, 13, 19) {real, imag} */,
  {32'h42edca6f, 32'hc22e1b4a} /* (29, 13, 18) {real, imag} */,
  {32'h4198163c, 32'hc154f7c5} /* (29, 13, 17) {real, imag} */,
  {32'hc2684b15, 32'h00000000} /* (29, 13, 16) {real, imag} */,
  {32'h4198163c, 32'h4154f7c5} /* (29, 13, 15) {real, imag} */,
  {32'h42edca6f, 32'h422e1b4a} /* (29, 13, 14) {real, imag} */,
  {32'hc26c3b6e, 32'h4244a7a4} /* (29, 13, 13) {real, imag} */,
  {32'hc1946cc1, 32'h414dfb98} /* (29, 13, 12) {real, imag} */,
  {32'h423a95e7, 32'hc27d31bc} /* (29, 13, 11) {real, imag} */,
  {32'h42768b20, 32'hc22573d9} /* (29, 13, 10) {real, imag} */,
  {32'hc2d76482, 32'hc2c24a86} /* (29, 13, 9) {real, imag} */,
  {32'hc127f05a, 32'h42d097a4} /* (29, 13, 8) {real, imag} */,
  {32'hc0b910cc, 32'hc1b1e822} /* (29, 13, 7) {real, imag} */,
  {32'h42e60748, 32'hc2e94ffe} /* (29, 13, 6) {real, imag} */,
  {32'h438cd8e1, 32'h431775b4} /* (29, 13, 5) {real, imag} */,
  {32'hc3531b27, 32'hc2ee22ec} /* (29, 13, 4) {real, imag} */,
  {32'hc242621c, 32'h420eb58f} /* (29, 13, 3) {real, imag} */,
  {32'h4474df0c, 32'h431d230a} /* (29, 13, 2) {real, imag} */,
  {32'hc4e1bee2, 32'hc32a7014} /* (29, 13, 1) {real, imag} */,
  {32'hc4c48d93, 32'h00000000} /* (29, 13, 0) {real, imag} */,
  {32'hc4c5a03d, 32'h42cac73c} /* (29, 12, 31) {real, imag} */,
  {32'h4438d5ee, 32'hc2685028} /* (29, 12, 30) {real, imag} */,
  {32'h3fcb95c0, 32'hc3038b7a} /* (29, 12, 29) {real, imag} */,
  {32'hc3692c0a, 32'h412f757c} /* (29, 12, 28) {real, imag} */,
  {32'h42e33637, 32'hc3b4fca4} /* (29, 12, 27) {real, imag} */,
  {32'hc2a9d120, 32'hc2c7a309} /* (29, 12, 26) {real, imag} */,
  {32'hc1f2bdc9, 32'hc07ceff0} /* (29, 12, 25) {real, imag} */,
  {32'hc18b6f11, 32'hc32d66a4} /* (29, 12, 24) {real, imag} */,
  {32'h4264f50d, 32'h428342e4} /* (29, 12, 23) {real, imag} */,
  {32'h436b550e, 32'h41994f44} /* (29, 12, 22) {real, imag} */,
  {32'h42338fbd, 32'hc2aa11c4} /* (29, 12, 21) {real, imag} */,
  {32'h421501be, 32'h413f134b} /* (29, 12, 20) {real, imag} */,
  {32'hc2835dde, 32'hc26279a5} /* (29, 12, 19) {real, imag} */,
  {32'h422ce591, 32'h41f763c3} /* (29, 12, 18) {real, imag} */,
  {32'h41cc9168, 32'h419f1cef} /* (29, 12, 17) {real, imag} */,
  {32'h4134d0e4, 32'h00000000} /* (29, 12, 16) {real, imag} */,
  {32'h41cc9168, 32'hc19f1cef} /* (29, 12, 15) {real, imag} */,
  {32'h422ce591, 32'hc1f763c3} /* (29, 12, 14) {real, imag} */,
  {32'hc2835dde, 32'h426279a5} /* (29, 12, 13) {real, imag} */,
  {32'h421501be, 32'hc13f134b} /* (29, 12, 12) {real, imag} */,
  {32'h42338fbd, 32'h42aa11c4} /* (29, 12, 11) {real, imag} */,
  {32'h436b550e, 32'hc1994f44} /* (29, 12, 10) {real, imag} */,
  {32'h4264f50d, 32'hc28342e4} /* (29, 12, 9) {real, imag} */,
  {32'hc18b6f11, 32'h432d66a4} /* (29, 12, 8) {real, imag} */,
  {32'hc1f2bdc9, 32'h407ceff0} /* (29, 12, 7) {real, imag} */,
  {32'hc2a9d120, 32'h42c7a309} /* (29, 12, 6) {real, imag} */,
  {32'h42e33637, 32'h43b4fca4} /* (29, 12, 5) {real, imag} */,
  {32'hc3692c0a, 32'hc12f757c} /* (29, 12, 4) {real, imag} */,
  {32'h3fcb95c0, 32'h43038b7a} /* (29, 12, 3) {real, imag} */,
  {32'h4438d5ee, 32'h42685028} /* (29, 12, 2) {real, imag} */,
  {32'hc4c5a03d, 32'hc2cac73c} /* (29, 12, 1) {real, imag} */,
  {32'hc4959e46, 32'h00000000} /* (29, 12, 0) {real, imag} */,
  {32'hc45c9a5b, 32'h425e8914} /* (29, 11, 31) {real, imag} */,
  {32'h43d67563, 32'hc1275f50} /* (29, 11, 30) {real, imag} */,
  {32'hc2ce521c, 32'hc2be18e8} /* (29, 11, 29) {real, imag} */,
  {32'hbfd27380, 32'hc29afcc7} /* (29, 11, 28) {real, imag} */,
  {32'h422f8fe0, 32'hc3ae5b63} /* (29, 11, 27) {real, imag} */,
  {32'hc2c5159d, 32'hc1915984} /* (29, 11, 26) {real, imag} */,
  {32'h42d2e654, 32'hc2368087} /* (29, 11, 25) {real, imag} */,
  {32'h42088f16, 32'h427f87df} /* (29, 11, 24) {real, imag} */,
  {32'h421c0556, 32'h42af06b1} /* (29, 11, 23) {real, imag} */,
  {32'h40bc310e, 32'h3f5a7ee0} /* (29, 11, 22) {real, imag} */,
  {32'hc2a6e4b6, 32'hc2c42a34} /* (29, 11, 21) {real, imag} */,
  {32'h40d46518, 32'hc26cd6ec} /* (29, 11, 20) {real, imag} */,
  {32'hbf44dbc0, 32'h42468b98} /* (29, 11, 19) {real, imag} */,
  {32'hc2bc4313, 32'hc23345d4} /* (29, 11, 18) {real, imag} */,
  {32'h40f48468, 32'h3f9ee9f0} /* (29, 11, 17) {real, imag} */,
  {32'h42725a7c, 32'h00000000} /* (29, 11, 16) {real, imag} */,
  {32'h40f48468, 32'hbf9ee9f0} /* (29, 11, 15) {real, imag} */,
  {32'hc2bc4313, 32'h423345d4} /* (29, 11, 14) {real, imag} */,
  {32'hbf44dbc0, 32'hc2468b98} /* (29, 11, 13) {real, imag} */,
  {32'h40d46518, 32'h426cd6ec} /* (29, 11, 12) {real, imag} */,
  {32'hc2a6e4b6, 32'h42c42a34} /* (29, 11, 11) {real, imag} */,
  {32'h40bc310e, 32'hbf5a7ee0} /* (29, 11, 10) {real, imag} */,
  {32'h421c0556, 32'hc2af06b1} /* (29, 11, 9) {real, imag} */,
  {32'h42088f16, 32'hc27f87df} /* (29, 11, 8) {real, imag} */,
  {32'h42d2e654, 32'h42368087} /* (29, 11, 7) {real, imag} */,
  {32'hc2c5159d, 32'h41915984} /* (29, 11, 6) {real, imag} */,
  {32'h422f8fe0, 32'h43ae5b63} /* (29, 11, 5) {real, imag} */,
  {32'hbfd27380, 32'h429afcc7} /* (29, 11, 4) {real, imag} */,
  {32'hc2ce521c, 32'h42be18e8} /* (29, 11, 3) {real, imag} */,
  {32'h43d67563, 32'h41275f50} /* (29, 11, 2) {real, imag} */,
  {32'hc45c9a5b, 32'hc25e8914} /* (29, 11, 1) {real, imag} */,
  {32'hc45e227c, 32'h00000000} /* (29, 11, 0) {real, imag} */,
  {32'h4417f932, 32'hc2be4df5} /* (29, 10, 31) {real, imag} */,
  {32'hc2465698, 32'h41137100} /* (29, 10, 30) {real, imag} */,
  {32'hc313365e, 32'h42bff9c5} /* (29, 10, 29) {real, imag} */,
  {32'h4212fb08, 32'hc2356436} /* (29, 10, 28) {real, imag} */,
  {32'hc27351b6, 32'hc17a8e4c} /* (29, 10, 27) {real, imag} */,
  {32'h4244b53f, 32'h404e57c0} /* (29, 10, 26) {real, imag} */,
  {32'h42ff0a73, 32'h426faaca} /* (29, 10, 25) {real, imag} */,
  {32'hc1b5af16, 32'hc20417e2} /* (29, 10, 24) {real, imag} */,
  {32'h41db93dd, 32'h418b30e2} /* (29, 10, 23) {real, imag} */,
  {32'hc2054f3f, 32'hc191e27d} /* (29, 10, 22) {real, imag} */,
  {32'hc30241d7, 32'h42c1a84c} /* (29, 10, 21) {real, imag} */,
  {32'h42ff75ac, 32'h41d13828} /* (29, 10, 20) {real, imag} */,
  {32'h408ada70, 32'hc0efa2e4} /* (29, 10, 19) {real, imag} */,
  {32'h42a0a9d1, 32'hc2f7e9f7} /* (29, 10, 18) {real, imag} */,
  {32'h41164b7a, 32'hc22d8e20} /* (29, 10, 17) {real, imag} */,
  {32'hc2133327, 32'h00000000} /* (29, 10, 16) {real, imag} */,
  {32'h41164b7a, 32'h422d8e20} /* (29, 10, 15) {real, imag} */,
  {32'h42a0a9d1, 32'h42f7e9f7} /* (29, 10, 14) {real, imag} */,
  {32'h408ada70, 32'h40efa2e4} /* (29, 10, 13) {real, imag} */,
  {32'h42ff75ac, 32'hc1d13828} /* (29, 10, 12) {real, imag} */,
  {32'hc30241d7, 32'hc2c1a84c} /* (29, 10, 11) {real, imag} */,
  {32'hc2054f3f, 32'h4191e27d} /* (29, 10, 10) {real, imag} */,
  {32'h41db93dd, 32'hc18b30e2} /* (29, 10, 9) {real, imag} */,
  {32'hc1b5af16, 32'h420417e2} /* (29, 10, 8) {real, imag} */,
  {32'h42ff0a73, 32'hc26faaca} /* (29, 10, 7) {real, imag} */,
  {32'h4244b53f, 32'hc04e57c0} /* (29, 10, 6) {real, imag} */,
  {32'hc27351b6, 32'h417a8e4c} /* (29, 10, 5) {real, imag} */,
  {32'h4212fb08, 32'h42356436} /* (29, 10, 4) {real, imag} */,
  {32'hc313365e, 32'hc2bff9c5} /* (29, 10, 3) {real, imag} */,
  {32'hc2465698, 32'hc1137100} /* (29, 10, 2) {real, imag} */,
  {32'h4417f932, 32'h42be4df5} /* (29, 10, 1) {real, imag} */,
  {32'h4298e2d0, 32'h00000000} /* (29, 10, 0) {real, imag} */,
  {32'h44b6cba4, 32'hc3780ca4} /* (29, 9, 31) {real, imag} */,
  {32'hc3dac215, 32'h4355f0ac} /* (29, 9, 30) {real, imag} */,
  {32'hc2e6199e, 32'hc1e07478} /* (29, 9, 29) {real, imag} */,
  {32'h421daca7, 32'hc2f772ae} /* (29, 9, 28) {real, imag} */,
  {32'hc36da061, 32'hc1b6d00c} /* (29, 9, 27) {real, imag} */,
  {32'hc3057635, 32'h41e9fb4e} /* (29, 9, 26) {real, imag} */,
  {32'h42e5a67c, 32'h4063b7b0} /* (29, 9, 25) {real, imag} */,
  {32'hc2938e4c, 32'h4185a42d} /* (29, 9, 24) {real, imag} */,
  {32'h42e78151, 32'hc2365637} /* (29, 9, 23) {real, imag} */,
  {32'h43185995, 32'h42d3c6e8} /* (29, 9, 22) {real, imag} */,
  {32'hc27393b0, 32'hc1363bb8} /* (29, 9, 21) {real, imag} */,
  {32'h428003e8, 32'h418751b0} /* (29, 9, 20) {real, imag} */,
  {32'hc14ced1e, 32'hc19d4ca8} /* (29, 9, 19) {real, imag} */,
  {32'h4185246e, 32'h4156de11} /* (29, 9, 18) {real, imag} */,
  {32'hc1884052, 32'h4267b48d} /* (29, 9, 17) {real, imag} */,
  {32'hc16cbd7c, 32'h00000000} /* (29, 9, 16) {real, imag} */,
  {32'hc1884052, 32'hc267b48d} /* (29, 9, 15) {real, imag} */,
  {32'h4185246e, 32'hc156de11} /* (29, 9, 14) {real, imag} */,
  {32'hc14ced1e, 32'h419d4ca8} /* (29, 9, 13) {real, imag} */,
  {32'h428003e8, 32'hc18751b0} /* (29, 9, 12) {real, imag} */,
  {32'hc27393b0, 32'h41363bb8} /* (29, 9, 11) {real, imag} */,
  {32'h43185995, 32'hc2d3c6e8} /* (29, 9, 10) {real, imag} */,
  {32'h42e78151, 32'h42365637} /* (29, 9, 9) {real, imag} */,
  {32'hc2938e4c, 32'hc185a42d} /* (29, 9, 8) {real, imag} */,
  {32'h42e5a67c, 32'hc063b7b0} /* (29, 9, 7) {real, imag} */,
  {32'hc3057635, 32'hc1e9fb4e} /* (29, 9, 6) {real, imag} */,
  {32'hc36da061, 32'h41b6d00c} /* (29, 9, 5) {real, imag} */,
  {32'h421daca7, 32'h42f772ae} /* (29, 9, 4) {real, imag} */,
  {32'hc2e6199e, 32'h41e07478} /* (29, 9, 3) {real, imag} */,
  {32'hc3dac215, 32'hc355f0ac} /* (29, 9, 2) {real, imag} */,
  {32'h44b6cba4, 32'h43780ca4} /* (29, 9, 1) {real, imag} */,
  {32'h440cf812, 32'h00000000} /* (29, 9, 0) {real, imag} */,
  {32'h44cf5a30, 32'hc3859354} /* (29, 8, 31) {real, imag} */,
  {32'hc3e9e048, 32'h43ec9c90} /* (29, 8, 30) {real, imag} */,
  {32'h413233ec, 32'h41b93c6e} /* (29, 8, 29) {real, imag} */,
  {32'h42ee2f76, 32'hc2d1f58f} /* (29, 8, 28) {real, imag} */,
  {32'hc3939ab0, 32'h40a97b78} /* (29, 8, 27) {real, imag} */,
  {32'h4137edbc, 32'hbf8a2b80} /* (29, 8, 26) {real, imag} */,
  {32'hc23fa0a4, 32'hc2e747c4} /* (29, 8, 25) {real, imag} */,
  {32'hc2609657, 32'h42889d01} /* (29, 8, 24) {real, imag} */,
  {32'hc2a6d594, 32'h42de58d1} /* (29, 8, 23) {real, imag} */,
  {32'h422690a5, 32'h41c7b4f8} /* (29, 8, 22) {real, imag} */,
  {32'h4182c7f6, 32'h42e2c866} /* (29, 8, 21) {real, imag} */,
  {32'hc20b5751, 32'hc13444dc} /* (29, 8, 20) {real, imag} */,
  {32'hc1cc2bab, 32'h4252802c} /* (29, 8, 19) {real, imag} */,
  {32'hc281180a, 32'hc20e4df2} /* (29, 8, 18) {real, imag} */,
  {32'hbf6b5b80, 32'hc296ee2e} /* (29, 8, 17) {real, imag} */,
  {32'hc019040e, 32'h00000000} /* (29, 8, 16) {real, imag} */,
  {32'hbf6b5b80, 32'h4296ee2e} /* (29, 8, 15) {real, imag} */,
  {32'hc281180a, 32'h420e4df2} /* (29, 8, 14) {real, imag} */,
  {32'hc1cc2bab, 32'hc252802c} /* (29, 8, 13) {real, imag} */,
  {32'hc20b5751, 32'h413444dc} /* (29, 8, 12) {real, imag} */,
  {32'h4182c7f6, 32'hc2e2c866} /* (29, 8, 11) {real, imag} */,
  {32'h422690a5, 32'hc1c7b4f8} /* (29, 8, 10) {real, imag} */,
  {32'hc2a6d594, 32'hc2de58d1} /* (29, 8, 9) {real, imag} */,
  {32'hc2609657, 32'hc2889d01} /* (29, 8, 8) {real, imag} */,
  {32'hc23fa0a4, 32'h42e747c4} /* (29, 8, 7) {real, imag} */,
  {32'h4137edbc, 32'h3f8a2b80} /* (29, 8, 6) {real, imag} */,
  {32'hc3939ab0, 32'hc0a97b78} /* (29, 8, 5) {real, imag} */,
  {32'h42ee2f76, 32'h42d1f58f} /* (29, 8, 4) {real, imag} */,
  {32'h413233ec, 32'hc1b93c6e} /* (29, 8, 3) {real, imag} */,
  {32'hc3e9e048, 32'hc3ec9c90} /* (29, 8, 2) {real, imag} */,
  {32'h44cf5a30, 32'h43859354} /* (29, 8, 1) {real, imag} */,
  {32'h4438ab54, 32'h00000000} /* (29, 8, 0) {real, imag} */,
  {32'h44ce65e8, 32'hc386c533} /* (29, 7, 31) {real, imag} */,
  {32'hc41c637c, 32'h43dd5147} /* (29, 7, 30) {real, imag} */,
  {32'h41ddcffe, 32'h4309917a} /* (29, 7, 29) {real, imag} */,
  {32'h427ea625, 32'hc206e6fc} /* (29, 7, 28) {real, imag} */,
  {32'hc3887c0a, 32'h42943a5a} /* (29, 7, 27) {real, imag} */,
  {32'h419a1292, 32'hc2df410a} /* (29, 7, 26) {real, imag} */,
  {32'hc307c5cc, 32'hc240baaf} /* (29, 7, 25) {real, imag} */,
  {32'hc1aa381a, 32'h428283f9} /* (29, 7, 24) {real, imag} */,
  {32'hc2a89a92, 32'h4250be5e} /* (29, 7, 23) {real, imag} */,
  {32'hc2c77785, 32'hc09b7a6c} /* (29, 7, 22) {real, imag} */,
  {32'h42c4c874, 32'h3ed5b200} /* (29, 7, 21) {real, imag} */,
  {32'hc1c0fdc4, 32'hc234e207} /* (29, 7, 20) {real, imag} */,
  {32'h427c984e, 32'h42b8f729} /* (29, 7, 19) {real, imag} */,
  {32'hc1cdf5d4, 32'hc0c263a3} /* (29, 7, 18) {real, imag} */,
  {32'h42041ded, 32'hc1cf45d4} /* (29, 7, 17) {real, imag} */,
  {32'h4236b301, 32'h00000000} /* (29, 7, 16) {real, imag} */,
  {32'h42041ded, 32'h41cf45d4} /* (29, 7, 15) {real, imag} */,
  {32'hc1cdf5d4, 32'h40c263a3} /* (29, 7, 14) {real, imag} */,
  {32'h427c984e, 32'hc2b8f729} /* (29, 7, 13) {real, imag} */,
  {32'hc1c0fdc4, 32'h4234e207} /* (29, 7, 12) {real, imag} */,
  {32'h42c4c874, 32'hbed5b200} /* (29, 7, 11) {real, imag} */,
  {32'hc2c77785, 32'h409b7a6c} /* (29, 7, 10) {real, imag} */,
  {32'hc2a89a92, 32'hc250be5e} /* (29, 7, 9) {real, imag} */,
  {32'hc1aa381a, 32'hc28283f9} /* (29, 7, 8) {real, imag} */,
  {32'hc307c5cc, 32'h4240baaf} /* (29, 7, 7) {real, imag} */,
  {32'h419a1292, 32'h42df410a} /* (29, 7, 6) {real, imag} */,
  {32'hc3887c0a, 32'hc2943a5a} /* (29, 7, 5) {real, imag} */,
  {32'h427ea625, 32'h4206e6fc} /* (29, 7, 4) {real, imag} */,
  {32'h41ddcffe, 32'hc309917a} /* (29, 7, 3) {real, imag} */,
  {32'hc41c637c, 32'hc3dd5147} /* (29, 7, 2) {real, imag} */,
  {32'h44ce65e8, 32'h4386c533} /* (29, 7, 1) {real, imag} */,
  {32'h44495449, 32'h00000000} /* (29, 7, 0) {real, imag} */,
  {32'h44c74bf7, 32'hc40713ce} /* (29, 6, 31) {real, imag} */,
  {32'hc3fdbe0a, 32'h440dd4af} /* (29, 6, 30) {real, imag} */,
  {32'h414e2724, 32'h415e6594} /* (29, 6, 29) {real, imag} */,
  {32'hbf8ed960, 32'hc2164e16} /* (29, 6, 28) {real, imag} */,
  {32'hc2ddcdd0, 32'hc1c1af04} /* (29, 6, 27) {real, imag} */,
  {32'hc28616ae, 32'hc290a6df} /* (29, 6, 26) {real, imag} */,
  {32'h4294d9a2, 32'hbf034ee0} /* (29, 6, 25) {real, imag} */,
  {32'hc2aca3e2, 32'h43132e3a} /* (29, 6, 24) {real, imag} */,
  {32'hc262cd45, 32'hbffc5be0} /* (29, 6, 23) {real, imag} */,
  {32'hc1bf53cc, 32'h4293779d} /* (29, 6, 22) {real, imag} */,
  {32'hc13ef64c, 32'h413e7620} /* (29, 6, 21) {real, imag} */,
  {32'hc22f9c34, 32'hc20640e6} /* (29, 6, 20) {real, imag} */,
  {32'h40adf2c2, 32'hc2975a3e} /* (29, 6, 19) {real, imag} */,
  {32'h4153edbf, 32'h42453856} /* (29, 6, 18) {real, imag} */,
  {32'hc1036896, 32'hc194413e} /* (29, 6, 17) {real, imag} */,
  {32'hc2974b17, 32'h00000000} /* (29, 6, 16) {real, imag} */,
  {32'hc1036896, 32'h4194413e} /* (29, 6, 15) {real, imag} */,
  {32'h4153edbf, 32'hc2453856} /* (29, 6, 14) {real, imag} */,
  {32'h40adf2c2, 32'h42975a3e} /* (29, 6, 13) {real, imag} */,
  {32'hc22f9c34, 32'h420640e6} /* (29, 6, 12) {real, imag} */,
  {32'hc13ef64c, 32'hc13e7620} /* (29, 6, 11) {real, imag} */,
  {32'hc1bf53cc, 32'hc293779d} /* (29, 6, 10) {real, imag} */,
  {32'hc262cd45, 32'h3ffc5be0} /* (29, 6, 9) {real, imag} */,
  {32'hc2aca3e2, 32'hc3132e3a} /* (29, 6, 8) {real, imag} */,
  {32'h4294d9a2, 32'h3f034ee0} /* (29, 6, 7) {real, imag} */,
  {32'hc28616ae, 32'h4290a6df} /* (29, 6, 6) {real, imag} */,
  {32'hc2ddcdd0, 32'h41c1af04} /* (29, 6, 5) {real, imag} */,
  {32'hbf8ed960, 32'h42164e16} /* (29, 6, 4) {real, imag} */,
  {32'h414e2724, 32'hc15e6594} /* (29, 6, 3) {real, imag} */,
  {32'hc3fdbe0a, 32'hc40dd4af} /* (29, 6, 2) {real, imag} */,
  {32'h44c74bf7, 32'h440713ce} /* (29, 6, 1) {real, imag} */,
  {32'h443d85ba, 32'h00000000} /* (29, 6, 0) {real, imag} */,
  {32'h449f0de9, 32'hc487b207} /* (29, 5, 31) {real, imag} */,
  {32'hc30f2fd4, 32'h445a93b9} /* (29, 5, 30) {real, imag} */,
  {32'hc22eefb6, 32'hc2205258} /* (29, 5, 29) {real, imag} */,
  {32'hc268a38e, 32'hc22865a4} /* (29, 5, 28) {real, imag} */,
  {32'hc321dda4, 32'h42a91dd4} /* (29, 5, 27) {real, imag} */,
  {32'hc19e6b56, 32'hc2974843} /* (29, 5, 26) {real, imag} */,
  {32'hc1eacfb0, 32'hc29f258e} /* (29, 5, 25) {real, imag} */,
  {32'h4210e8da, 32'h4333572a} /* (29, 5, 24) {real, imag} */,
  {32'h420819ce, 32'h41b7ea91} /* (29, 5, 23) {real, imag} */,
  {32'h422e9d76, 32'h42ea0515} /* (29, 5, 22) {real, imag} */,
  {32'hc2986632, 32'h428776d0} /* (29, 5, 21) {real, imag} */,
  {32'hc0c30cc1, 32'hc0d67da0} /* (29, 5, 20) {real, imag} */,
  {32'h41bfac90, 32'hc2926e98} /* (29, 5, 19) {real, imag} */,
  {32'hc18aaf10, 32'h42a6bbe9} /* (29, 5, 18) {real, imag} */,
  {32'hc11d2ac2, 32'hc2b54b1f} /* (29, 5, 17) {real, imag} */,
  {32'h426a9a6a, 32'h00000000} /* (29, 5, 16) {real, imag} */,
  {32'hc11d2ac2, 32'h42b54b1f} /* (29, 5, 15) {real, imag} */,
  {32'hc18aaf10, 32'hc2a6bbe9} /* (29, 5, 14) {real, imag} */,
  {32'h41bfac90, 32'h42926e98} /* (29, 5, 13) {real, imag} */,
  {32'hc0c30cc1, 32'h40d67da0} /* (29, 5, 12) {real, imag} */,
  {32'hc2986632, 32'hc28776d0} /* (29, 5, 11) {real, imag} */,
  {32'h422e9d76, 32'hc2ea0515} /* (29, 5, 10) {real, imag} */,
  {32'h420819ce, 32'hc1b7ea91} /* (29, 5, 9) {real, imag} */,
  {32'h4210e8da, 32'hc333572a} /* (29, 5, 8) {real, imag} */,
  {32'hc1eacfb0, 32'h429f258e} /* (29, 5, 7) {real, imag} */,
  {32'hc19e6b56, 32'h42974843} /* (29, 5, 6) {real, imag} */,
  {32'hc321dda4, 32'hc2a91dd4} /* (29, 5, 5) {real, imag} */,
  {32'hc268a38e, 32'h422865a4} /* (29, 5, 4) {real, imag} */,
  {32'hc22eefb6, 32'h42205258} /* (29, 5, 3) {real, imag} */,
  {32'hc30f2fd4, 32'hc45a93b9} /* (29, 5, 2) {real, imag} */,
  {32'h449f0de9, 32'h4487b207} /* (29, 5, 1) {real, imag} */,
  {32'h446f288e, 32'h00000000} /* (29, 5, 0) {real, imag} */,
  {32'h44573440, 32'hc4a54443} /* (29, 4, 31) {real, imag} */,
  {32'h4313c2fa, 32'h446ec296} /* (29, 4, 30) {real, imag} */,
  {32'hc2cfc438, 32'hc2be323e} /* (29, 4, 29) {real, imag} */,
  {32'hc36d5216, 32'h433d0ef1} /* (29, 4, 28) {real, imag} */,
  {32'hc28dedd0, 32'h41e86c32} /* (29, 4, 27) {real, imag} */,
  {32'hc239ec44, 32'hc15cad26} /* (29, 4, 26) {real, imag} */,
  {32'hc120f054, 32'hc2beb622} /* (29, 4, 25) {real, imag} */,
  {32'h4312e682, 32'h42e559c4} /* (29, 4, 24) {real, imag} */,
  {32'hc27d7809, 32'hc1e70467} /* (29, 4, 23) {real, imag} */,
  {32'hc24311d4, 32'h41e2ff79} /* (29, 4, 22) {real, imag} */,
  {32'h42336cfe, 32'hc2429a93} /* (29, 4, 21) {real, imag} */,
  {32'hc28ac309, 32'hc2536118} /* (29, 4, 20) {real, imag} */,
  {32'hc21277e9, 32'h3fc07480} /* (29, 4, 19) {real, imag} */,
  {32'h42619b3c, 32'hc29ab4b3} /* (29, 4, 18) {real, imag} */,
  {32'hc09b2309, 32'hc186b576} /* (29, 4, 17) {real, imag} */,
  {32'h427a0373, 32'h00000000} /* (29, 4, 16) {real, imag} */,
  {32'hc09b2309, 32'h4186b576} /* (29, 4, 15) {real, imag} */,
  {32'h42619b3c, 32'h429ab4b3} /* (29, 4, 14) {real, imag} */,
  {32'hc21277e9, 32'hbfc07480} /* (29, 4, 13) {real, imag} */,
  {32'hc28ac309, 32'h42536118} /* (29, 4, 12) {real, imag} */,
  {32'h42336cfe, 32'h42429a93} /* (29, 4, 11) {real, imag} */,
  {32'hc24311d4, 32'hc1e2ff79} /* (29, 4, 10) {real, imag} */,
  {32'hc27d7809, 32'h41e70467} /* (29, 4, 9) {real, imag} */,
  {32'h4312e682, 32'hc2e559c4} /* (29, 4, 8) {real, imag} */,
  {32'hc120f054, 32'h42beb622} /* (29, 4, 7) {real, imag} */,
  {32'hc239ec44, 32'h415cad26} /* (29, 4, 6) {real, imag} */,
  {32'hc28dedd0, 32'hc1e86c32} /* (29, 4, 5) {real, imag} */,
  {32'hc36d5216, 32'hc33d0ef1} /* (29, 4, 4) {real, imag} */,
  {32'hc2cfc438, 32'h42be323e} /* (29, 4, 3) {real, imag} */,
  {32'h4313c2fa, 32'hc46ec296} /* (29, 4, 2) {real, imag} */,
  {32'h44573440, 32'h44a54443} /* (29, 4, 1) {real, imag} */,
  {32'h44563e5f, 32'h00000000} /* (29, 4, 0) {real, imag} */,
  {32'h44124b7d, 32'hc4ab91be} /* (29, 3, 31) {real, imag} */,
  {32'h439c16e7, 32'h443b3ce8} /* (29, 3, 30) {real, imag} */,
  {32'hc31372d2, 32'hc2ea62d9} /* (29, 3, 29) {real, imag} */,
  {32'hc30c5b6b, 32'h4354ffdd} /* (29, 3, 28) {real, imag} */,
  {32'hc2d4f13c, 32'hc23cdb86} /* (29, 3, 27) {real, imag} */,
  {32'hc289fd74, 32'h41d2ec1a} /* (29, 3, 26) {real, imag} */,
  {32'hc20a3708, 32'hc2ddebff} /* (29, 3, 25) {real, imag} */,
  {32'h42782408, 32'h420a26c2} /* (29, 3, 24) {real, imag} */,
  {32'hc187a258, 32'h40b3f850} /* (29, 3, 23) {real, imag} */,
  {32'hc008f890, 32'h412357ec} /* (29, 3, 22) {real, imag} */,
  {32'h429cd9ea, 32'h428cdd34} /* (29, 3, 21) {real, imag} */,
  {32'hc14bc350, 32'hc251f9e8} /* (29, 3, 20) {real, imag} */,
  {32'h429aae67, 32'hc1b4a864} /* (29, 3, 19) {real, imag} */,
  {32'h413e7696, 32'hc21aab48} /* (29, 3, 18) {real, imag} */,
  {32'h40e5377e, 32'h41710080} /* (29, 3, 17) {real, imag} */,
  {32'h4196013e, 32'h00000000} /* (29, 3, 16) {real, imag} */,
  {32'h40e5377e, 32'hc1710080} /* (29, 3, 15) {real, imag} */,
  {32'h413e7696, 32'h421aab48} /* (29, 3, 14) {real, imag} */,
  {32'h429aae67, 32'h41b4a864} /* (29, 3, 13) {real, imag} */,
  {32'hc14bc350, 32'h4251f9e8} /* (29, 3, 12) {real, imag} */,
  {32'h429cd9ea, 32'hc28cdd34} /* (29, 3, 11) {real, imag} */,
  {32'hc008f890, 32'hc12357ec} /* (29, 3, 10) {real, imag} */,
  {32'hc187a258, 32'hc0b3f850} /* (29, 3, 9) {real, imag} */,
  {32'h42782408, 32'hc20a26c2} /* (29, 3, 8) {real, imag} */,
  {32'hc20a3708, 32'h42ddebff} /* (29, 3, 7) {real, imag} */,
  {32'hc289fd74, 32'hc1d2ec1a} /* (29, 3, 6) {real, imag} */,
  {32'hc2d4f13c, 32'h423cdb86} /* (29, 3, 5) {real, imag} */,
  {32'hc30c5b6b, 32'hc354ffdd} /* (29, 3, 4) {real, imag} */,
  {32'hc31372d2, 32'h42ea62d9} /* (29, 3, 3) {real, imag} */,
  {32'h439c16e7, 32'hc43b3ce8} /* (29, 3, 2) {real, imag} */,
  {32'h44124b7d, 32'h44ab91be} /* (29, 3, 1) {real, imag} */,
  {32'h4405d4d0, 32'h00000000} /* (29, 3, 0) {real, imag} */,
  {32'h440419d1, 32'hc4c10672} /* (29, 2, 31) {real, imag} */,
  {32'h43b392d4, 32'h441a253a} /* (29, 2, 30) {real, imag} */,
  {32'hc257c5c2, 32'hc2acea4a} /* (29, 2, 29) {real, imag} */,
  {32'hc29b7680, 32'h41c925e8} /* (29, 2, 28) {real, imag} */,
  {32'hc329306f, 32'hc2b2b84b} /* (29, 2, 27) {real, imag} */,
  {32'hc22404f3, 32'hbe2e0800} /* (29, 2, 26) {real, imag} */,
  {32'hc26c7aa5, 32'hc343c39a} /* (29, 2, 25) {real, imag} */,
  {32'h4222c19a, 32'h42832c82} /* (29, 2, 24) {real, imag} */,
  {32'h42cf7874, 32'h42717388} /* (29, 2, 23) {real, imag} */,
  {32'hc2380816, 32'h4223454e} /* (29, 2, 22) {real, imag} */,
  {32'hc1d779dc, 32'h41d10745} /* (29, 2, 21) {real, imag} */,
  {32'hc2b23b8f, 32'h4256749e} /* (29, 2, 20) {real, imag} */,
  {32'h421e5708, 32'h410a7d74} /* (29, 2, 19) {real, imag} */,
  {32'hc2159988, 32'h41068504} /* (29, 2, 18) {real, imag} */,
  {32'h42346dae, 32'h4184298b} /* (29, 2, 17) {real, imag} */,
  {32'hc1d45f0e, 32'h00000000} /* (29, 2, 16) {real, imag} */,
  {32'h42346dae, 32'hc184298b} /* (29, 2, 15) {real, imag} */,
  {32'hc2159988, 32'hc1068504} /* (29, 2, 14) {real, imag} */,
  {32'h421e5708, 32'hc10a7d74} /* (29, 2, 13) {real, imag} */,
  {32'hc2b23b8f, 32'hc256749e} /* (29, 2, 12) {real, imag} */,
  {32'hc1d779dc, 32'hc1d10745} /* (29, 2, 11) {real, imag} */,
  {32'hc2380816, 32'hc223454e} /* (29, 2, 10) {real, imag} */,
  {32'h42cf7874, 32'hc2717388} /* (29, 2, 9) {real, imag} */,
  {32'h4222c19a, 32'hc2832c82} /* (29, 2, 8) {real, imag} */,
  {32'hc26c7aa5, 32'h4343c39a} /* (29, 2, 7) {real, imag} */,
  {32'hc22404f3, 32'h3e2e0800} /* (29, 2, 6) {real, imag} */,
  {32'hc329306f, 32'h42b2b84b} /* (29, 2, 5) {real, imag} */,
  {32'hc29b7680, 32'hc1c925e8} /* (29, 2, 4) {real, imag} */,
  {32'hc257c5c2, 32'h42acea4a} /* (29, 2, 3) {real, imag} */,
  {32'h43b392d4, 32'hc41a253a} /* (29, 2, 2) {real, imag} */,
  {32'h440419d1, 32'h44c10672} /* (29, 2, 1) {real, imag} */,
  {32'h44138b47, 32'h00000000} /* (29, 2, 0) {real, imag} */,
  {32'h441234e4, 32'hc4ba2d6a} /* (29, 1, 31) {real, imag} */,
  {32'h432b0236, 32'h444f74c8} /* (29, 1, 30) {real, imag} */,
  {32'hc2eeaf3c, 32'hc1c4da00} /* (29, 1, 29) {real, imag} */,
  {32'hc14639c8, 32'h43515804} /* (29, 1, 28) {real, imag} */,
  {32'hc35d3e6d, 32'hc0ca86a4} /* (29, 1, 27) {real, imag} */,
  {32'hc27586a8, 32'hc128f706} /* (29, 1, 26) {real, imag} */,
  {32'h40bc3ee4, 32'hc2c504a2} /* (29, 1, 25) {real, imag} */,
  {32'h41bb55d0, 32'h420a18b6} /* (29, 1, 24) {real, imag} */,
  {32'h411b40fb, 32'hc2fd6545} /* (29, 1, 23) {real, imag} */,
  {32'h41615976, 32'h4209bb94} /* (29, 1, 22) {real, imag} */,
  {32'hc235f841, 32'h4141f784} /* (29, 1, 21) {real, imag} */,
  {32'hc202de0c, 32'hc266132a} /* (29, 1, 20) {real, imag} */,
  {32'h418d4537, 32'h421c9cbe} /* (29, 1, 19) {real, imag} */,
  {32'hc22eba58, 32'h4206b5dd} /* (29, 1, 18) {real, imag} */,
  {32'h4146fb1e, 32'h41ac45d2} /* (29, 1, 17) {real, imag} */,
  {32'h41ebf630, 32'h00000000} /* (29, 1, 16) {real, imag} */,
  {32'h4146fb1e, 32'hc1ac45d2} /* (29, 1, 15) {real, imag} */,
  {32'hc22eba58, 32'hc206b5dd} /* (29, 1, 14) {real, imag} */,
  {32'h418d4537, 32'hc21c9cbe} /* (29, 1, 13) {real, imag} */,
  {32'hc202de0c, 32'h4266132a} /* (29, 1, 12) {real, imag} */,
  {32'hc235f841, 32'hc141f784} /* (29, 1, 11) {real, imag} */,
  {32'h41615976, 32'hc209bb94} /* (29, 1, 10) {real, imag} */,
  {32'h411b40fb, 32'h42fd6545} /* (29, 1, 9) {real, imag} */,
  {32'h41bb55d0, 32'hc20a18b6} /* (29, 1, 8) {real, imag} */,
  {32'h40bc3ee4, 32'h42c504a2} /* (29, 1, 7) {real, imag} */,
  {32'hc27586a8, 32'h4128f706} /* (29, 1, 6) {real, imag} */,
  {32'hc35d3e6d, 32'h40ca86a4} /* (29, 1, 5) {real, imag} */,
  {32'hc14639c8, 32'hc3515804} /* (29, 1, 4) {real, imag} */,
  {32'hc2eeaf3c, 32'h41c4da00} /* (29, 1, 3) {real, imag} */,
  {32'h432b0236, 32'hc44f74c8} /* (29, 1, 2) {real, imag} */,
  {32'h441234e4, 32'h44ba2d6a} /* (29, 1, 1) {real, imag} */,
  {32'h44178606, 32'h00000000} /* (29, 1, 0) {real, imag} */,
  {32'h4419a5fe, 32'hc47400e8} /* (29, 0, 31) {real, imag} */,
  {32'hc1277780, 32'h44356381} /* (29, 0, 30) {real, imag} */,
  {32'hc2aa0c03, 32'hc217d734} /* (29, 0, 29) {real, imag} */,
  {32'h41c618c6, 32'h43268a50} /* (29, 0, 28) {real, imag} */,
  {32'hc3603c91, 32'hc23122e1} /* (29, 0, 27) {real, imag} */,
  {32'hc208921e, 32'hc175c1b0} /* (29, 0, 26) {real, imag} */,
  {32'hc1ed9c25, 32'h4187d9a1} /* (29, 0, 25) {real, imag} */,
  {32'hc1695899, 32'h41e4369b} /* (29, 0, 24) {real, imag} */,
  {32'h41263f42, 32'h41dc6545} /* (29, 0, 23) {real, imag} */,
  {32'hc2bbab87, 32'h4243c606} /* (29, 0, 22) {real, imag} */,
  {32'h42133345, 32'hc278b0e2} /* (29, 0, 21) {real, imag} */,
  {32'h41c04872, 32'hc25b5933} /* (29, 0, 20) {real, imag} */,
  {32'h4298dd8c, 32'h41950579} /* (29, 0, 19) {real, imag} */,
  {32'h42401740, 32'h41bc0b2d} /* (29, 0, 18) {real, imag} */,
  {32'hc1ff4dc0, 32'hc1332040} /* (29, 0, 17) {real, imag} */,
  {32'h4064ccd8, 32'h00000000} /* (29, 0, 16) {real, imag} */,
  {32'hc1ff4dc0, 32'h41332040} /* (29, 0, 15) {real, imag} */,
  {32'h42401740, 32'hc1bc0b2d} /* (29, 0, 14) {real, imag} */,
  {32'h4298dd8c, 32'hc1950579} /* (29, 0, 13) {real, imag} */,
  {32'h41c04872, 32'h425b5933} /* (29, 0, 12) {real, imag} */,
  {32'h42133345, 32'h4278b0e2} /* (29, 0, 11) {real, imag} */,
  {32'hc2bbab87, 32'hc243c606} /* (29, 0, 10) {real, imag} */,
  {32'h41263f42, 32'hc1dc6545} /* (29, 0, 9) {real, imag} */,
  {32'hc1695899, 32'hc1e4369b} /* (29, 0, 8) {real, imag} */,
  {32'hc1ed9c25, 32'hc187d9a1} /* (29, 0, 7) {real, imag} */,
  {32'hc208921e, 32'h4175c1b0} /* (29, 0, 6) {real, imag} */,
  {32'hc3603c91, 32'h423122e1} /* (29, 0, 5) {real, imag} */,
  {32'h41c618c6, 32'hc3268a50} /* (29, 0, 4) {real, imag} */,
  {32'hc2aa0c03, 32'h4217d734} /* (29, 0, 3) {real, imag} */,
  {32'hc1277780, 32'hc4356381} /* (29, 0, 2) {real, imag} */,
  {32'h4419a5fe, 32'h447400e8} /* (29, 0, 1) {real, imag} */,
  {32'h43cdc3cc, 32'h00000000} /* (29, 0, 0) {real, imag} */,
  {32'h44365d3a, 32'hc3d04c52} /* (28, 31, 31) {real, imag} */,
  {32'hc3ed51db, 32'h43ff2a52} /* (28, 31, 30) {real, imag} */,
  {32'hc2e344e0, 32'h40a517b4} /* (28, 31, 29) {real, imag} */,
  {32'h426dc76f, 32'h4348ef09} /* (28, 31, 28) {real, imag} */,
  {32'hc3006a4f, 32'h42d86c26} /* (28, 31, 27) {real, imag} */,
  {32'h41d01ff7, 32'hc16f4618} /* (28, 31, 26) {real, imag} */,
  {32'h41bd2b9a, 32'hc2165512} /* (28, 31, 25) {real, imag} */,
  {32'hc230b255, 32'hc15702a4} /* (28, 31, 24) {real, imag} */,
  {32'h4147ec46, 32'h427284db} /* (28, 31, 23) {real, imag} */,
  {32'hc1424d2c, 32'h40d62734} /* (28, 31, 22) {real, imag} */,
  {32'hc2310634, 32'hc100ae6a} /* (28, 31, 21) {real, imag} */,
  {32'hc1b7a544, 32'hc2396a37} /* (28, 31, 20) {real, imag} */,
  {32'hc285b1f6, 32'hc20801f3} /* (28, 31, 19) {real, imag} */,
  {32'h41388db2, 32'hc186a1d0} /* (28, 31, 18) {real, imag} */,
  {32'hc04128ec, 32'h41202cb8} /* (28, 31, 17) {real, imag} */,
  {32'h410c0fca, 32'h00000000} /* (28, 31, 16) {real, imag} */,
  {32'hc04128ec, 32'hc1202cb8} /* (28, 31, 15) {real, imag} */,
  {32'h41388db2, 32'h4186a1d0} /* (28, 31, 14) {real, imag} */,
  {32'hc285b1f6, 32'h420801f3} /* (28, 31, 13) {real, imag} */,
  {32'hc1b7a544, 32'h42396a37} /* (28, 31, 12) {real, imag} */,
  {32'hc2310634, 32'h4100ae6a} /* (28, 31, 11) {real, imag} */,
  {32'hc1424d2c, 32'hc0d62734} /* (28, 31, 10) {real, imag} */,
  {32'h4147ec46, 32'hc27284db} /* (28, 31, 9) {real, imag} */,
  {32'hc230b255, 32'h415702a4} /* (28, 31, 8) {real, imag} */,
  {32'h41bd2b9a, 32'h42165512} /* (28, 31, 7) {real, imag} */,
  {32'h41d01ff7, 32'h416f4618} /* (28, 31, 6) {real, imag} */,
  {32'hc3006a4f, 32'hc2d86c26} /* (28, 31, 5) {real, imag} */,
  {32'h426dc76f, 32'hc348ef09} /* (28, 31, 4) {real, imag} */,
  {32'hc2e344e0, 32'hc0a517b4} /* (28, 31, 3) {real, imag} */,
  {32'hc3ed51db, 32'hc3ff2a52} /* (28, 31, 2) {real, imag} */,
  {32'h44365d3a, 32'h43d04c52} /* (28, 31, 1) {real, imag} */,
  {32'h42e55e54, 32'h00000000} /* (28, 31, 0) {real, imag} */,
  {32'h44970e2d, 32'hc3751170} /* (28, 30, 31) {real, imag} */,
  {32'hc471707f, 32'h43eb0c90} /* (28, 30, 30) {real, imag} */,
  {32'hc30154de, 32'h416e37d0} /* (28, 30, 29) {real, imag} */,
  {32'h42e7afda, 32'h42e3e924} /* (28, 30, 28) {real, imag} */,
  {32'hc329f685, 32'h43159042} /* (28, 30, 27) {real, imag} */,
  {32'hc212c3a4, 32'hc2f489c0} /* (28, 30, 26) {real, imag} */,
  {32'h42a747a1, 32'hc28b2e10} /* (28, 30, 25) {real, imag} */,
  {32'h41aa7eb4, 32'hc28c4eec} /* (28, 30, 24) {real, imag} */,
  {32'hc2158316, 32'hc1ca23c8} /* (28, 30, 23) {real, imag} */,
  {32'h424c84a2, 32'hc1de2418} /* (28, 30, 22) {real, imag} */,
  {32'hc27214d0, 32'h42a7e5f9} /* (28, 30, 21) {real, imag} */,
  {32'hc211d6d7, 32'hc21021c0} /* (28, 30, 20) {real, imag} */,
  {32'hc2787619, 32'hc235b981} /* (28, 30, 19) {real, imag} */,
  {32'h41f1d281, 32'hc1c06b03} /* (28, 30, 18) {real, imag} */,
  {32'h4062c900, 32'h420bf806} /* (28, 30, 17) {real, imag} */,
  {32'hc2ae478b, 32'h00000000} /* (28, 30, 16) {real, imag} */,
  {32'h4062c900, 32'hc20bf806} /* (28, 30, 15) {real, imag} */,
  {32'h41f1d281, 32'h41c06b03} /* (28, 30, 14) {real, imag} */,
  {32'hc2787619, 32'h4235b981} /* (28, 30, 13) {real, imag} */,
  {32'hc211d6d7, 32'h421021c0} /* (28, 30, 12) {real, imag} */,
  {32'hc27214d0, 32'hc2a7e5f9} /* (28, 30, 11) {real, imag} */,
  {32'h424c84a2, 32'h41de2418} /* (28, 30, 10) {real, imag} */,
  {32'hc2158316, 32'h41ca23c8} /* (28, 30, 9) {real, imag} */,
  {32'h41aa7eb4, 32'h428c4eec} /* (28, 30, 8) {real, imag} */,
  {32'h42a747a1, 32'h428b2e10} /* (28, 30, 7) {real, imag} */,
  {32'hc212c3a4, 32'h42f489c0} /* (28, 30, 6) {real, imag} */,
  {32'hc329f685, 32'hc3159042} /* (28, 30, 5) {real, imag} */,
  {32'h42e7afda, 32'hc2e3e924} /* (28, 30, 4) {real, imag} */,
  {32'hc30154de, 32'hc16e37d0} /* (28, 30, 3) {real, imag} */,
  {32'hc471707f, 32'hc3eb0c90} /* (28, 30, 2) {real, imag} */,
  {32'h44970e2d, 32'h43751170} /* (28, 30, 1) {real, imag} */,
  {32'h438abf02, 32'h00000000} /* (28, 30, 0) {real, imag} */,
  {32'h44bace3e, 32'hc295bae8} /* (28, 29, 31) {real, imag} */,
  {32'hc482b72c, 32'h438116ed} /* (28, 29, 30) {real, imag} */,
  {32'hc3159429, 32'h41ceff40} /* (28, 29, 29) {real, imag} */,
  {32'h4305689a, 32'h4116ec80} /* (28, 29, 28) {real, imag} */,
  {32'hc3699dde, 32'h414dc170} /* (28, 29, 27) {real, imag} */,
  {32'h409da244, 32'hc0d54790} /* (28, 29, 26) {real, imag} */,
  {32'hc1f50dc4, 32'hc25bcbb0} /* (28, 29, 25) {real, imag} */,
  {32'hc250ce82, 32'h421e8fc9} /* (28, 29, 24) {real, imag} */,
  {32'h42d546cb, 32'hc24c2ed6} /* (28, 29, 23) {real, imag} */,
  {32'h41b80fda, 32'hc2a7d6c7} /* (28, 29, 22) {real, imag} */,
  {32'hc2929944, 32'h4037b300} /* (28, 29, 21) {real, imag} */,
  {32'hc2c4aaa2, 32'hc22029ea} /* (28, 29, 20) {real, imag} */,
  {32'h4223aa9c, 32'h42740d03} /* (28, 29, 19) {real, imag} */,
  {32'hbf4ee1c0, 32'hc179ef3e} /* (28, 29, 18) {real, imag} */,
  {32'h422d971b, 32'h410845de} /* (28, 29, 17) {real, imag} */,
  {32'hc12b3414, 32'h00000000} /* (28, 29, 16) {real, imag} */,
  {32'h422d971b, 32'hc10845de} /* (28, 29, 15) {real, imag} */,
  {32'hbf4ee1c0, 32'h4179ef3e} /* (28, 29, 14) {real, imag} */,
  {32'h4223aa9c, 32'hc2740d03} /* (28, 29, 13) {real, imag} */,
  {32'hc2c4aaa2, 32'h422029ea} /* (28, 29, 12) {real, imag} */,
  {32'hc2929944, 32'hc037b300} /* (28, 29, 11) {real, imag} */,
  {32'h41b80fda, 32'h42a7d6c7} /* (28, 29, 10) {real, imag} */,
  {32'h42d546cb, 32'h424c2ed6} /* (28, 29, 9) {real, imag} */,
  {32'hc250ce82, 32'hc21e8fc9} /* (28, 29, 8) {real, imag} */,
  {32'hc1f50dc4, 32'h425bcbb0} /* (28, 29, 7) {real, imag} */,
  {32'h409da244, 32'h40d54790} /* (28, 29, 6) {real, imag} */,
  {32'hc3699dde, 32'hc14dc170} /* (28, 29, 5) {real, imag} */,
  {32'h4305689a, 32'hc116ec80} /* (28, 29, 4) {real, imag} */,
  {32'hc3159429, 32'hc1ceff40} /* (28, 29, 3) {real, imag} */,
  {32'hc482b72c, 32'hc38116ed} /* (28, 29, 2) {real, imag} */,
  {32'h44bace3e, 32'h4295bae8} /* (28, 29, 1) {real, imag} */,
  {32'h43649846, 32'h00000000} /* (28, 29, 0) {real, imag} */,
  {32'h44bd3a62, 32'h42ad5c70} /* (28, 28, 31) {real, imag} */,
  {32'hc49992ce, 32'h43875e6e} /* (28, 28, 30) {real, imag} */,
  {32'hc20ad1cf, 32'hc1b38dab} /* (28, 28, 29) {real, imag} */,
  {32'h43113822, 32'hc212c5dd} /* (28, 28, 28) {real, imag} */,
  {32'hc3bcc3a6, 32'h431b1a43} /* (28, 28, 27) {real, imag} */,
  {32'h41c67a8f, 32'hc22c89c6} /* (28, 28, 26) {real, imag} */,
  {32'h4189c07c, 32'hc2fcb1ab} /* (28, 28, 25) {real, imag} */,
  {32'hc274a0a9, 32'h42b9f786} /* (28, 28, 24) {real, imag} */,
  {32'h42785214, 32'hc24578c6} /* (28, 28, 23) {real, imag} */,
  {32'h41ee89ba, 32'hc2a6b48c} /* (28, 28, 22) {real, imag} */,
  {32'hc1696f60, 32'h4289276f} /* (28, 28, 21) {real, imag} */,
  {32'hc1ff94a5, 32'hc2dd5d4c} /* (28, 28, 20) {real, imag} */,
  {32'hc245e0be, 32'h4277b96a} /* (28, 28, 19) {real, imag} */,
  {32'hc121c348, 32'hc2204c2c} /* (28, 28, 18) {real, imag} */,
  {32'h41900398, 32'h41f615e0} /* (28, 28, 17) {real, imag} */,
  {32'h42db37de, 32'h00000000} /* (28, 28, 16) {real, imag} */,
  {32'h41900398, 32'hc1f615e0} /* (28, 28, 15) {real, imag} */,
  {32'hc121c348, 32'h42204c2c} /* (28, 28, 14) {real, imag} */,
  {32'hc245e0be, 32'hc277b96a} /* (28, 28, 13) {real, imag} */,
  {32'hc1ff94a5, 32'h42dd5d4c} /* (28, 28, 12) {real, imag} */,
  {32'hc1696f60, 32'hc289276f} /* (28, 28, 11) {real, imag} */,
  {32'h41ee89ba, 32'h42a6b48c} /* (28, 28, 10) {real, imag} */,
  {32'h42785214, 32'h424578c6} /* (28, 28, 9) {real, imag} */,
  {32'hc274a0a9, 32'hc2b9f786} /* (28, 28, 8) {real, imag} */,
  {32'h4189c07c, 32'h42fcb1ab} /* (28, 28, 7) {real, imag} */,
  {32'h41c67a8f, 32'h422c89c6} /* (28, 28, 6) {real, imag} */,
  {32'hc3bcc3a6, 32'hc31b1a43} /* (28, 28, 5) {real, imag} */,
  {32'h43113822, 32'h4212c5dd} /* (28, 28, 4) {real, imag} */,
  {32'hc20ad1cf, 32'h41b38dab} /* (28, 28, 3) {real, imag} */,
  {32'hc49992ce, 32'hc3875e6e} /* (28, 28, 2) {real, imag} */,
  {32'h44bd3a62, 32'hc2ad5c70} /* (28, 28, 1) {real, imag} */,
  {32'h43e008e2, 32'h00000000} /* (28, 28, 0) {real, imag} */,
  {32'h44b65eea, 32'h4337d9b4} /* (28, 27, 31) {real, imag} */,
  {32'hc491c7cc, 32'h4396959a} /* (28, 27, 30) {real, imag} */,
  {32'hc1664230, 32'hc33e2028} /* (28, 27, 29) {real, imag} */,
  {32'h42858894, 32'hc3051ef8} /* (28, 27, 28) {real, imag} */,
  {32'hc3810036, 32'h433e6510} /* (28, 27, 27) {real, imag} */,
  {32'hc20f5cfd, 32'hc1760ba8} /* (28, 27, 26) {real, imag} */,
  {32'h418ffcd2, 32'hbf3db280} /* (28, 27, 25) {real, imag} */,
  {32'hc264692e, 32'h43230d8c} /* (28, 27, 24) {real, imag} */,
  {32'h42841df4, 32'hc1bf6d7e} /* (28, 27, 23) {real, imag} */,
  {32'hc22d19f8, 32'hc1c545a8} /* (28, 27, 22) {real, imag} */,
  {32'hc281d7c4, 32'h42200be0} /* (28, 27, 21) {real, imag} */,
  {32'hc13ced18, 32'hc2917de4} /* (28, 27, 20) {real, imag} */,
  {32'h4294d56c, 32'hc311a7f0} /* (28, 27, 19) {real, imag} */,
  {32'h412b18f0, 32'h423ffa5c} /* (28, 27, 18) {real, imag} */,
  {32'h4278c4ae, 32'h42a0fad3} /* (28, 27, 17) {real, imag} */,
  {32'hc2b99a08, 32'h00000000} /* (28, 27, 16) {real, imag} */,
  {32'h4278c4ae, 32'hc2a0fad3} /* (28, 27, 15) {real, imag} */,
  {32'h412b18f0, 32'hc23ffa5c} /* (28, 27, 14) {real, imag} */,
  {32'h4294d56c, 32'h4311a7f0} /* (28, 27, 13) {real, imag} */,
  {32'hc13ced18, 32'h42917de4} /* (28, 27, 12) {real, imag} */,
  {32'hc281d7c4, 32'hc2200be0} /* (28, 27, 11) {real, imag} */,
  {32'hc22d19f8, 32'h41c545a8} /* (28, 27, 10) {real, imag} */,
  {32'h42841df4, 32'h41bf6d7e} /* (28, 27, 9) {real, imag} */,
  {32'hc264692e, 32'hc3230d8c} /* (28, 27, 8) {real, imag} */,
  {32'h418ffcd2, 32'h3f3db280} /* (28, 27, 7) {real, imag} */,
  {32'hc20f5cfd, 32'h41760ba8} /* (28, 27, 6) {real, imag} */,
  {32'hc3810036, 32'hc33e6510} /* (28, 27, 5) {real, imag} */,
  {32'h42858894, 32'h43051ef8} /* (28, 27, 4) {real, imag} */,
  {32'hc1664230, 32'h433e2028} /* (28, 27, 3) {real, imag} */,
  {32'hc491c7cc, 32'hc396959a} /* (28, 27, 2) {real, imag} */,
  {32'h44b65eea, 32'hc337d9b4} /* (28, 27, 1) {real, imag} */,
  {32'h441befb2, 32'h00000000} /* (28, 27, 0) {real, imag} */,
  {32'h44b1e26b, 32'h42c7159c} /* (28, 26, 31) {real, imag} */,
  {32'hc495b62c, 32'h437096b4} /* (28, 26, 30) {real, imag} */,
  {32'h4296bfd2, 32'hc23aad6a} /* (28, 26, 29) {real, imag} */,
  {32'h433a51be, 32'hc2ca576c} /* (28, 26, 28) {real, imag} */,
  {32'hc2b4361e, 32'h4345a722} /* (28, 26, 27) {real, imag} */,
  {32'hc133e4a4, 32'hc2307a98} /* (28, 26, 26) {real, imag} */,
  {32'h42ad4a9e, 32'hc2f2b5d8} /* (28, 26, 25) {real, imag} */,
  {32'h413b33f9, 32'h429416db} /* (28, 26, 24) {real, imag} */,
  {32'hc1bdc854, 32'h42a1b72f} /* (28, 26, 23) {real, imag} */,
  {32'hc2bc9289, 32'hc1ad6290} /* (28, 26, 22) {real, imag} */,
  {32'h424d30bc, 32'h3f5e5b5c} /* (28, 26, 21) {real, imag} */,
  {32'h4252512e, 32'h42441af4} /* (28, 26, 20) {real, imag} */,
  {32'hbf5b42c0, 32'hc218dcd1} /* (28, 26, 19) {real, imag} */,
  {32'hc2cd8b90, 32'h42db74d8} /* (28, 26, 18) {real, imag} */,
  {32'h424028a6, 32'hc211363a} /* (28, 26, 17) {real, imag} */,
  {32'h40219908, 32'h00000000} /* (28, 26, 16) {real, imag} */,
  {32'h424028a6, 32'h4211363a} /* (28, 26, 15) {real, imag} */,
  {32'hc2cd8b90, 32'hc2db74d8} /* (28, 26, 14) {real, imag} */,
  {32'hbf5b42c0, 32'h4218dcd1} /* (28, 26, 13) {real, imag} */,
  {32'h4252512e, 32'hc2441af4} /* (28, 26, 12) {real, imag} */,
  {32'h424d30bc, 32'hbf5e5b5c} /* (28, 26, 11) {real, imag} */,
  {32'hc2bc9289, 32'h41ad6290} /* (28, 26, 10) {real, imag} */,
  {32'hc1bdc854, 32'hc2a1b72f} /* (28, 26, 9) {real, imag} */,
  {32'h413b33f9, 32'hc29416db} /* (28, 26, 8) {real, imag} */,
  {32'h42ad4a9e, 32'h42f2b5d8} /* (28, 26, 7) {real, imag} */,
  {32'hc133e4a4, 32'h42307a98} /* (28, 26, 6) {real, imag} */,
  {32'hc2b4361e, 32'hc345a722} /* (28, 26, 5) {real, imag} */,
  {32'h433a51be, 32'h42ca576c} /* (28, 26, 4) {real, imag} */,
  {32'h4296bfd2, 32'h423aad6a} /* (28, 26, 3) {real, imag} */,
  {32'hc495b62c, 32'hc37096b4} /* (28, 26, 2) {real, imag} */,
  {32'h44b1e26b, 32'hc2c7159c} /* (28, 26, 1) {real, imag} */,
  {32'h43cdc814, 32'h00000000} /* (28, 26, 0) {real, imag} */,
  {32'h44a11918, 32'hc1155c90} /* (28, 25, 31) {real, imag} */,
  {32'hc48a0f34, 32'h4377453c} /* (28, 25, 30) {real, imag} */,
  {32'h419ec148, 32'hc26cf162} /* (28, 25, 29) {real, imag} */,
  {32'h4357f94d, 32'hc31c07f3} /* (28, 25, 28) {real, imag} */,
  {32'hc3058dcf, 32'h418cacf8} /* (28, 25, 27) {real, imag} */,
  {32'h4258d20d, 32'hc1ef2507} /* (28, 25, 26) {real, imag} */,
  {32'h42fd9b3a, 32'hc2d9d300} /* (28, 25, 25) {real, imag} */,
  {32'hc20cd180, 32'h420bff98} /* (28, 25, 24) {real, imag} */,
  {32'hc0c33eb8, 32'h42ab2cc0} /* (28, 25, 23) {real, imag} */,
  {32'hc1884dbc, 32'hc20ea075} /* (28, 25, 22) {real, imag} */,
  {32'hc2b55acd, 32'hc2d01700} /* (28, 25, 21) {real, imag} */,
  {32'h4286cbba, 32'h40e3700c} /* (28, 25, 20) {real, imag} */,
  {32'h420172ec, 32'h414d3bc8} /* (28, 25, 19) {real, imag} */,
  {32'hbf0a0e80, 32'h41d4e0fd} /* (28, 25, 18) {real, imag} */,
  {32'hbff319f0, 32'hc1822a96} /* (28, 25, 17) {real, imag} */,
  {32'hc1d31e6b, 32'h00000000} /* (28, 25, 16) {real, imag} */,
  {32'hbff319f0, 32'h41822a96} /* (28, 25, 15) {real, imag} */,
  {32'hbf0a0e80, 32'hc1d4e0fd} /* (28, 25, 14) {real, imag} */,
  {32'h420172ec, 32'hc14d3bc8} /* (28, 25, 13) {real, imag} */,
  {32'h4286cbba, 32'hc0e3700c} /* (28, 25, 12) {real, imag} */,
  {32'hc2b55acd, 32'h42d01700} /* (28, 25, 11) {real, imag} */,
  {32'hc1884dbc, 32'h420ea075} /* (28, 25, 10) {real, imag} */,
  {32'hc0c33eb8, 32'hc2ab2cc0} /* (28, 25, 9) {real, imag} */,
  {32'hc20cd180, 32'hc20bff98} /* (28, 25, 8) {real, imag} */,
  {32'h42fd9b3a, 32'h42d9d300} /* (28, 25, 7) {real, imag} */,
  {32'h4258d20d, 32'h41ef2507} /* (28, 25, 6) {real, imag} */,
  {32'hc3058dcf, 32'hc18cacf8} /* (28, 25, 5) {real, imag} */,
  {32'h4357f94d, 32'h431c07f3} /* (28, 25, 4) {real, imag} */,
  {32'h419ec148, 32'h426cf162} /* (28, 25, 3) {real, imag} */,
  {32'hc48a0f34, 32'hc377453c} /* (28, 25, 2) {real, imag} */,
  {32'h44a11918, 32'h41155c90} /* (28, 25, 1) {real, imag} */,
  {32'h441bcfa3, 32'h00000000} /* (28, 25, 0) {real, imag} */,
  {32'h44a1267c, 32'hc21e6ece} /* (28, 24, 31) {real, imag} */,
  {32'hc499d6ca, 32'h43a73b18} /* (28, 24, 30) {real, imag} */,
  {32'hc1c98e88, 32'hc3403452} /* (28, 24, 29) {real, imag} */,
  {32'h434d3346, 32'h42526b68} /* (28, 24, 28) {real, imag} */,
  {32'hc2940552, 32'h415dcdf0} /* (28, 24, 27) {real, imag} */,
  {32'hc1e62f41, 32'h42b6a532} /* (28, 24, 26) {real, imag} */,
  {32'hc26bbdda, 32'hc316963b} /* (28, 24, 25) {real, imag} */,
  {32'h427c8ca0, 32'h427ad9ce} /* (28, 24, 24) {real, imag} */,
  {32'hc2b10b73, 32'h421a82aa} /* (28, 24, 23) {real, imag} */,
  {32'hc1992642, 32'h41b5fe28} /* (28, 24, 22) {real, imag} */,
  {32'hc242792e, 32'h4287cbbb} /* (28, 24, 21) {real, imag} */,
  {32'h4112cd5c, 32'h41cbd66a} /* (28, 24, 20) {real, imag} */,
  {32'h42c2244d, 32'h42925f98} /* (28, 24, 19) {real, imag} */,
  {32'h40ea06d8, 32'hc1c46e59} /* (28, 24, 18) {real, imag} */,
  {32'hc1b17048, 32'hc2863064} /* (28, 24, 17) {real, imag} */,
  {32'hc192978b, 32'h00000000} /* (28, 24, 16) {real, imag} */,
  {32'hc1b17048, 32'h42863064} /* (28, 24, 15) {real, imag} */,
  {32'h40ea06d8, 32'h41c46e59} /* (28, 24, 14) {real, imag} */,
  {32'h42c2244d, 32'hc2925f98} /* (28, 24, 13) {real, imag} */,
  {32'h4112cd5c, 32'hc1cbd66a} /* (28, 24, 12) {real, imag} */,
  {32'hc242792e, 32'hc287cbbb} /* (28, 24, 11) {real, imag} */,
  {32'hc1992642, 32'hc1b5fe28} /* (28, 24, 10) {real, imag} */,
  {32'hc2b10b73, 32'hc21a82aa} /* (28, 24, 9) {real, imag} */,
  {32'h427c8ca0, 32'hc27ad9ce} /* (28, 24, 8) {real, imag} */,
  {32'hc26bbdda, 32'h4316963b} /* (28, 24, 7) {real, imag} */,
  {32'hc1e62f41, 32'hc2b6a532} /* (28, 24, 6) {real, imag} */,
  {32'hc2940552, 32'hc15dcdf0} /* (28, 24, 5) {real, imag} */,
  {32'h434d3346, 32'hc2526b68} /* (28, 24, 4) {real, imag} */,
  {32'hc1c98e88, 32'h43403452} /* (28, 24, 3) {real, imag} */,
  {32'hc499d6ca, 32'hc3a73b18} /* (28, 24, 2) {real, imag} */,
  {32'h44a1267c, 32'h421e6ece} /* (28, 24, 1) {real, imag} */,
  {32'h4432906c, 32'h00000000} /* (28, 24, 0) {real, imag} */,
  {32'h4485969e, 32'hc2d5239a} /* (28, 23, 31) {real, imag} */,
  {32'hc477d9f6, 32'h43147a4f} /* (28, 23, 30) {real, imag} */,
  {32'hc1910422, 32'hc2c3737f} /* (28, 23, 29) {real, imag} */,
  {32'h42b34655, 32'hc2586a78} /* (28, 23, 28) {real, imag} */,
  {32'hc23bf354, 32'h4343817a} /* (28, 23, 27) {real, imag} */,
  {32'h40237770, 32'h42347ef6} /* (28, 23, 26) {real, imag} */,
  {32'hc26bdece, 32'hc33f38e4} /* (28, 23, 25) {real, imag} */,
  {32'hc1f6f299, 32'h42defbf8} /* (28, 23, 24) {real, imag} */,
  {32'hc2c4c674, 32'hc28370ab} /* (28, 23, 23) {real, imag} */,
  {32'hc19ebadc, 32'h4221708c} /* (28, 23, 22) {real, imag} */,
  {32'h42a061b3, 32'h424c22cb} /* (28, 23, 21) {real, imag} */,
  {32'h41fced74, 32'hc25ee2dc} /* (28, 23, 20) {real, imag} */,
  {32'hc223a1e2, 32'hc1c0c748} /* (28, 23, 19) {real, imag} */,
  {32'h4182f90e, 32'h428008cb} /* (28, 23, 18) {real, imag} */,
  {32'h42341ba9, 32'h426c9759} /* (28, 23, 17) {real, imag} */,
  {32'hc2d30014, 32'h00000000} /* (28, 23, 16) {real, imag} */,
  {32'h42341ba9, 32'hc26c9759} /* (28, 23, 15) {real, imag} */,
  {32'h4182f90e, 32'hc28008cb} /* (28, 23, 14) {real, imag} */,
  {32'hc223a1e2, 32'h41c0c748} /* (28, 23, 13) {real, imag} */,
  {32'h41fced74, 32'h425ee2dc} /* (28, 23, 12) {real, imag} */,
  {32'h42a061b3, 32'hc24c22cb} /* (28, 23, 11) {real, imag} */,
  {32'hc19ebadc, 32'hc221708c} /* (28, 23, 10) {real, imag} */,
  {32'hc2c4c674, 32'h428370ab} /* (28, 23, 9) {real, imag} */,
  {32'hc1f6f299, 32'hc2defbf8} /* (28, 23, 8) {real, imag} */,
  {32'hc26bdece, 32'h433f38e4} /* (28, 23, 7) {real, imag} */,
  {32'h40237770, 32'hc2347ef6} /* (28, 23, 6) {real, imag} */,
  {32'hc23bf354, 32'hc343817a} /* (28, 23, 5) {real, imag} */,
  {32'h42b34655, 32'h42586a78} /* (28, 23, 4) {real, imag} */,
  {32'hc1910422, 32'h42c3737f} /* (28, 23, 3) {real, imag} */,
  {32'hc477d9f6, 32'hc3147a4f} /* (28, 23, 2) {real, imag} */,
  {32'h4485969e, 32'h42d5239a} /* (28, 23, 1) {real, imag} */,
  {32'h443b063a, 32'h00000000} /* (28, 23, 0) {real, imag} */,
  {32'h44295648, 32'hc0639fa0} /* (28, 22, 31) {real, imag} */,
  {32'hc3eb1098, 32'h420393c5} /* (28, 22, 30) {real, imag} */,
  {32'h42212e5a, 32'hc2cd7a91} /* (28, 22, 29) {real, imag} */,
  {32'hc0eecf90, 32'hc2cf0af8} /* (28, 22, 28) {real, imag} */,
  {32'hc3145658, 32'h41ffb712} /* (28, 22, 27) {real, imag} */,
  {32'hc291d2cc, 32'h42292486} /* (28, 22, 26) {real, imag} */,
  {32'hc1f5261a, 32'hc3166c28} /* (28, 22, 25) {real, imag} */,
  {32'hc26c96e6, 32'h41977f02} /* (28, 22, 24) {real, imag} */,
  {32'hc1ab6fb7, 32'h429148ce} /* (28, 22, 23) {real, imag} */,
  {32'hc169504e, 32'h42aedba7} /* (28, 22, 22) {real, imag} */,
  {32'h4205a3b0, 32'h42720685} /* (28, 22, 21) {real, imag} */,
  {32'hc19f8c8c, 32'h429fc474} /* (28, 22, 20) {real, imag} */,
  {32'h41fa46b5, 32'hc01c2640} /* (28, 22, 19) {real, imag} */,
  {32'hc1effe33, 32'h4191b284} /* (28, 22, 18) {real, imag} */,
  {32'h41af401c, 32'h40907248} /* (28, 22, 17) {real, imag} */,
  {32'h41e21ee4, 32'h00000000} /* (28, 22, 16) {real, imag} */,
  {32'h41af401c, 32'hc0907248} /* (28, 22, 15) {real, imag} */,
  {32'hc1effe33, 32'hc191b284} /* (28, 22, 14) {real, imag} */,
  {32'h41fa46b5, 32'h401c2640} /* (28, 22, 13) {real, imag} */,
  {32'hc19f8c8c, 32'hc29fc474} /* (28, 22, 12) {real, imag} */,
  {32'h4205a3b0, 32'hc2720685} /* (28, 22, 11) {real, imag} */,
  {32'hc169504e, 32'hc2aedba7} /* (28, 22, 10) {real, imag} */,
  {32'hc1ab6fb7, 32'hc29148ce} /* (28, 22, 9) {real, imag} */,
  {32'hc26c96e6, 32'hc1977f02} /* (28, 22, 8) {real, imag} */,
  {32'hc1f5261a, 32'h43166c28} /* (28, 22, 7) {real, imag} */,
  {32'hc291d2cc, 32'hc2292486} /* (28, 22, 6) {real, imag} */,
  {32'hc3145658, 32'hc1ffb712} /* (28, 22, 5) {real, imag} */,
  {32'hc0eecf90, 32'h42cf0af8} /* (28, 22, 4) {real, imag} */,
  {32'h42212e5a, 32'h42cd7a91} /* (28, 22, 3) {real, imag} */,
  {32'hc3eb1098, 32'hc20393c5} /* (28, 22, 2) {real, imag} */,
  {32'h44295648, 32'h40639fa0} /* (28, 22, 1) {real, imag} */,
  {32'h44246f99, 32'h00000000} /* (28, 22, 0) {real, imag} */,
  {32'hc2c6581c, 32'h42001a94} /* (28, 21, 31) {real, imag} */,
  {32'hc1e6fbe8, 32'h4133f540} /* (28, 21, 30) {real, imag} */,
  {32'h425ad882, 32'hc1c4b74c} /* (28, 21, 29) {real, imag} */,
  {32'hc2388ff4, 32'hc0849ae8} /* (28, 21, 28) {real, imag} */,
  {32'hc256c3ff, 32'hc20ee0e7} /* (28, 21, 27) {real, imag} */,
  {32'hc262593d, 32'h4218fc2a} /* (28, 21, 26) {real, imag} */,
  {32'h42583076, 32'h422bb030} /* (28, 21, 25) {real, imag} */,
  {32'h42a5a0ca, 32'h42b4c6f9} /* (28, 21, 24) {real, imag} */,
  {32'h4213526c, 32'hc2235060} /* (28, 21, 23) {real, imag} */,
  {32'h425fa561, 32'h425481ab} /* (28, 21, 22) {real, imag} */,
  {32'hc1cba790, 32'h42d9e1f0} /* (28, 21, 21) {real, imag} */,
  {32'hc1bd4b2c, 32'hc260c016} /* (28, 21, 20) {real, imag} */,
  {32'hc1a8772c, 32'hc0c8dba0} /* (28, 21, 19) {real, imag} */,
  {32'hc2ca9278, 32'hc2141690} /* (28, 21, 18) {real, imag} */,
  {32'hbf3ee9c0, 32'hc2408030} /* (28, 21, 17) {real, imag} */,
  {32'hc0aea170, 32'h00000000} /* (28, 21, 16) {real, imag} */,
  {32'hbf3ee9c0, 32'h42408030} /* (28, 21, 15) {real, imag} */,
  {32'hc2ca9278, 32'h42141690} /* (28, 21, 14) {real, imag} */,
  {32'hc1a8772c, 32'h40c8dba0} /* (28, 21, 13) {real, imag} */,
  {32'hc1bd4b2c, 32'h4260c016} /* (28, 21, 12) {real, imag} */,
  {32'hc1cba790, 32'hc2d9e1f0} /* (28, 21, 11) {real, imag} */,
  {32'h425fa561, 32'hc25481ab} /* (28, 21, 10) {real, imag} */,
  {32'h4213526c, 32'h42235060} /* (28, 21, 9) {real, imag} */,
  {32'h42a5a0ca, 32'hc2b4c6f9} /* (28, 21, 8) {real, imag} */,
  {32'h42583076, 32'hc22bb030} /* (28, 21, 7) {real, imag} */,
  {32'hc262593d, 32'hc218fc2a} /* (28, 21, 6) {real, imag} */,
  {32'hc256c3ff, 32'h420ee0e7} /* (28, 21, 5) {real, imag} */,
  {32'hc2388ff4, 32'h40849ae8} /* (28, 21, 4) {real, imag} */,
  {32'h425ad882, 32'h41c4b74c} /* (28, 21, 3) {real, imag} */,
  {32'hc1e6fbe8, 32'hc133f540} /* (28, 21, 2) {real, imag} */,
  {32'hc2c6581c, 32'hc2001a94} /* (28, 21, 1) {real, imag} */,
  {32'hbef32c00, 32'h00000000} /* (28, 21, 0) {real, imag} */,
  {32'hc492d9e6, 32'h43663e28} /* (28, 20, 31) {real, imag} */,
  {32'h4404c0a6, 32'hc34948c5} /* (28, 20, 30) {real, imag} */,
  {32'h4322e8d9, 32'hc2b0fa18} /* (28, 20, 29) {real, imag} */,
  {32'hc339610a, 32'h41f7beac} /* (28, 20, 28) {real, imag} */,
  {32'h42c2c111, 32'hc1dbfda8} /* (28, 20, 27) {real, imag} */,
  {32'h420c139c, 32'hc2460f26} /* (28, 20, 26) {real, imag} */,
  {32'h42099e0d, 32'h422a5907} /* (28, 20, 25) {real, imag} */,
  {32'h41437336, 32'hc2e34c18} /* (28, 20, 24) {real, imag} */,
  {32'h427c6ef8, 32'hc27f7b30} /* (28, 20, 23) {real, imag} */,
  {32'h4334135b, 32'h4237d0de} /* (28, 20, 22) {real, imag} */,
  {32'h431980e9, 32'h42761046} /* (28, 20, 21) {real, imag} */,
  {32'h41abacea, 32'h3ff6d280} /* (28, 20, 20) {real, imag} */,
  {32'hc23d1232, 32'h41926321} /* (28, 20, 19) {real, imag} */,
  {32'h42035434, 32'hbfe3ab00} /* (28, 20, 18) {real, imag} */,
  {32'h412ec2c0, 32'h427bb2c8} /* (28, 20, 17) {real, imag} */,
  {32'hc28056c5, 32'h00000000} /* (28, 20, 16) {real, imag} */,
  {32'h412ec2c0, 32'hc27bb2c8} /* (28, 20, 15) {real, imag} */,
  {32'h42035434, 32'h3fe3ab00} /* (28, 20, 14) {real, imag} */,
  {32'hc23d1232, 32'hc1926321} /* (28, 20, 13) {real, imag} */,
  {32'h41abacea, 32'hbff6d280} /* (28, 20, 12) {real, imag} */,
  {32'h431980e9, 32'hc2761046} /* (28, 20, 11) {real, imag} */,
  {32'h4334135b, 32'hc237d0de} /* (28, 20, 10) {real, imag} */,
  {32'h427c6ef8, 32'h427f7b30} /* (28, 20, 9) {real, imag} */,
  {32'h41437336, 32'h42e34c18} /* (28, 20, 8) {real, imag} */,
  {32'h42099e0d, 32'hc22a5907} /* (28, 20, 7) {real, imag} */,
  {32'h420c139c, 32'h42460f26} /* (28, 20, 6) {real, imag} */,
  {32'h42c2c111, 32'h41dbfda8} /* (28, 20, 5) {real, imag} */,
  {32'hc339610a, 32'hc1f7beac} /* (28, 20, 4) {real, imag} */,
  {32'h4322e8d9, 32'h42b0fa18} /* (28, 20, 3) {real, imag} */,
  {32'h4404c0a6, 32'h434948c5} /* (28, 20, 2) {real, imag} */,
  {32'hc492d9e6, 32'hc3663e28} /* (28, 20, 1) {real, imag} */,
  {32'hc422adfe, 32'h00000000} /* (28, 20, 0) {real, imag} */,
  {32'hc4cd16d2, 32'h4386ce36} /* (28, 19, 31) {real, imag} */,
  {32'h4429588d, 32'hc3698e90} /* (28, 19, 30) {real, imag} */,
  {32'h41969f38, 32'hc2ea2df8} /* (28, 19, 29) {real, imag} */,
  {32'hc2fb0b68, 32'h41f42046} /* (28, 19, 28) {real, imag} */,
  {32'h428d395a, 32'h41c24978} /* (28, 19, 27) {real, imag} */,
  {32'hc28a9825, 32'hc23ccd73} /* (28, 19, 26) {real, imag} */,
  {32'hc25f188e, 32'h422fece0} /* (28, 19, 25) {real, imag} */,
  {32'hc132fc00, 32'hc2dd023c} /* (28, 19, 24) {real, imag} */,
  {32'h4256b3ec, 32'hc0f7c826} /* (28, 19, 23) {real, imag} */,
  {32'h42c5b552, 32'hc10c007c} /* (28, 19, 22) {real, imag} */,
  {32'hc203bc13, 32'hc02e8058} /* (28, 19, 21) {real, imag} */,
  {32'hc1610fe8, 32'h3fab3c64} /* (28, 19, 20) {real, imag} */,
  {32'hc26c7eeb, 32'hc0af3568} /* (28, 19, 19) {real, imag} */,
  {32'hc28eb912, 32'hc22e01dc} /* (28, 19, 18) {real, imag} */,
  {32'hc22b69f5, 32'hc20b2866} /* (28, 19, 17) {real, imag} */,
  {32'hc261f6dc, 32'h00000000} /* (28, 19, 16) {real, imag} */,
  {32'hc22b69f5, 32'h420b2866} /* (28, 19, 15) {real, imag} */,
  {32'hc28eb912, 32'h422e01dc} /* (28, 19, 14) {real, imag} */,
  {32'hc26c7eeb, 32'h40af3568} /* (28, 19, 13) {real, imag} */,
  {32'hc1610fe8, 32'hbfab3c64} /* (28, 19, 12) {real, imag} */,
  {32'hc203bc13, 32'h402e8058} /* (28, 19, 11) {real, imag} */,
  {32'h42c5b552, 32'h410c007c} /* (28, 19, 10) {real, imag} */,
  {32'h4256b3ec, 32'h40f7c826} /* (28, 19, 9) {real, imag} */,
  {32'hc132fc00, 32'h42dd023c} /* (28, 19, 8) {real, imag} */,
  {32'hc25f188e, 32'hc22fece0} /* (28, 19, 7) {real, imag} */,
  {32'hc28a9825, 32'h423ccd73} /* (28, 19, 6) {real, imag} */,
  {32'h428d395a, 32'hc1c24978} /* (28, 19, 5) {real, imag} */,
  {32'hc2fb0b68, 32'hc1f42046} /* (28, 19, 4) {real, imag} */,
  {32'h41969f38, 32'h42ea2df8} /* (28, 19, 3) {real, imag} */,
  {32'h4429588d, 32'h43698e90} /* (28, 19, 2) {real, imag} */,
  {32'hc4cd16d2, 32'hc386ce36} /* (28, 19, 1) {real, imag} */,
  {32'hc48e4cc6, 32'h00000000} /* (28, 19, 0) {real, imag} */,
  {32'hc4e9aaab, 32'h43c240e8} /* (28, 18, 31) {real, imag} */,
  {32'h4463df0b, 32'hc3ac505a} /* (28, 18, 30) {real, imag} */,
  {32'hc281bb72, 32'hc0a08d60} /* (28, 18, 29) {real, imag} */,
  {32'hc28edc86, 32'h430c81a8} /* (28, 18, 28) {real, imag} */,
  {32'h43474709, 32'hc2eda588} /* (28, 18, 27) {real, imag} */,
  {32'hc2fd11f6, 32'hc20183b7} /* (28, 18, 26) {real, imag} */,
  {32'h41c00045, 32'h42b41c7e} /* (28, 18, 25) {real, imag} */,
  {32'h4252fa6b, 32'hc2c36303} /* (28, 18, 24) {real, imag} */,
  {32'h40b23128, 32'hc2df202e} /* (28, 18, 23) {real, imag} */,
  {32'h428d588a, 32'h40f85298} /* (28, 18, 22) {real, imag} */,
  {32'hc1c6fb08, 32'h41221130} /* (28, 18, 21) {real, imag} */,
  {32'hc0ebab40, 32'hc214924e} /* (28, 18, 20) {real, imag} */,
  {32'hc294fbeb, 32'h4278ef70} /* (28, 18, 19) {real, imag} */,
  {32'hc1c6d14b, 32'hc25822ae} /* (28, 18, 18) {real, imag} */,
  {32'hc2988a7b, 32'h423091fa} /* (28, 18, 17) {real, imag} */,
  {32'hc0feba91, 32'h00000000} /* (28, 18, 16) {real, imag} */,
  {32'hc2988a7b, 32'hc23091fa} /* (28, 18, 15) {real, imag} */,
  {32'hc1c6d14b, 32'h425822ae} /* (28, 18, 14) {real, imag} */,
  {32'hc294fbeb, 32'hc278ef70} /* (28, 18, 13) {real, imag} */,
  {32'hc0ebab40, 32'h4214924e} /* (28, 18, 12) {real, imag} */,
  {32'hc1c6fb08, 32'hc1221130} /* (28, 18, 11) {real, imag} */,
  {32'h428d588a, 32'hc0f85298} /* (28, 18, 10) {real, imag} */,
  {32'h40b23128, 32'h42df202e} /* (28, 18, 9) {real, imag} */,
  {32'h4252fa6b, 32'h42c36303} /* (28, 18, 8) {real, imag} */,
  {32'h41c00045, 32'hc2b41c7e} /* (28, 18, 7) {real, imag} */,
  {32'hc2fd11f6, 32'h420183b7} /* (28, 18, 6) {real, imag} */,
  {32'h43474709, 32'h42eda588} /* (28, 18, 5) {real, imag} */,
  {32'hc28edc86, 32'hc30c81a8} /* (28, 18, 4) {real, imag} */,
  {32'hc281bb72, 32'h40a08d60} /* (28, 18, 3) {real, imag} */,
  {32'h4463df0b, 32'h43ac505a} /* (28, 18, 2) {real, imag} */,
  {32'hc4e9aaab, 32'hc3c240e8} /* (28, 18, 1) {real, imag} */,
  {32'hc4b7e1c5, 32'h00000000} /* (28, 18, 0) {real, imag} */,
  {32'hc4f27d43, 32'h43f8d990} /* (28, 17, 31) {real, imag} */,
  {32'h4473e612, 32'hc345f708} /* (28, 17, 30) {real, imag} */,
  {32'h42cc1a0c, 32'hc250e180} /* (28, 17, 29) {real, imag} */,
  {32'hc2a071c5, 32'h42c92f48} /* (28, 17, 28) {real, imag} */,
  {32'h43412984, 32'hc23004a2} /* (28, 17, 27) {real, imag} */,
  {32'h418bb190, 32'hc216c8a1} /* (28, 17, 26) {real, imag} */,
  {32'h42dd42c4, 32'h42846666} /* (28, 17, 25) {real, imag} */,
  {32'h423fff44, 32'hbfce0a90} /* (28, 17, 24) {real, imag} */,
  {32'h41bde91e, 32'hc1b7f5ca} /* (28, 17, 23) {real, imag} */,
  {32'hc2f8020f, 32'hc2a5e3d0} /* (28, 17, 22) {real, imag} */,
  {32'hc1ecf772, 32'hc21c1408} /* (28, 17, 21) {real, imag} */,
  {32'h411f148a, 32'h411bf754} /* (28, 17, 20) {real, imag} */,
  {32'h41d363de, 32'hc280f300} /* (28, 17, 19) {real, imag} */,
  {32'h41ce3728, 32'h3f80af00} /* (28, 17, 18) {real, imag} */,
  {32'hc220e2a5, 32'h4267a770} /* (28, 17, 17) {real, imag} */,
  {32'h431fff0e, 32'h00000000} /* (28, 17, 16) {real, imag} */,
  {32'hc220e2a5, 32'hc267a770} /* (28, 17, 15) {real, imag} */,
  {32'h41ce3728, 32'hbf80af00} /* (28, 17, 14) {real, imag} */,
  {32'h41d363de, 32'h4280f300} /* (28, 17, 13) {real, imag} */,
  {32'h411f148a, 32'hc11bf754} /* (28, 17, 12) {real, imag} */,
  {32'hc1ecf772, 32'h421c1408} /* (28, 17, 11) {real, imag} */,
  {32'hc2f8020f, 32'h42a5e3d0} /* (28, 17, 10) {real, imag} */,
  {32'h41bde91e, 32'h41b7f5ca} /* (28, 17, 9) {real, imag} */,
  {32'h423fff44, 32'h3fce0a90} /* (28, 17, 8) {real, imag} */,
  {32'h42dd42c4, 32'hc2846666} /* (28, 17, 7) {real, imag} */,
  {32'h418bb190, 32'h4216c8a1} /* (28, 17, 6) {real, imag} */,
  {32'h43412984, 32'h423004a2} /* (28, 17, 5) {real, imag} */,
  {32'hc2a071c5, 32'hc2c92f48} /* (28, 17, 4) {real, imag} */,
  {32'h42cc1a0c, 32'h4250e180} /* (28, 17, 3) {real, imag} */,
  {32'h4473e612, 32'h4345f708} /* (28, 17, 2) {real, imag} */,
  {32'hc4f27d43, 32'hc3f8d990} /* (28, 17, 1) {real, imag} */,
  {32'hc4d094f4, 32'h00000000} /* (28, 17, 0) {real, imag} */,
  {32'hc4f21890, 32'h43afb89e} /* (28, 16, 31) {real, imag} */,
  {32'h447ecd50, 32'hc345907a} /* (28, 16, 30) {real, imag} */,
  {32'h428e49e5, 32'h4198ffd6} /* (28, 16, 29) {real, imag} */,
  {32'hc2a7a401, 32'h4320d283} /* (28, 16, 28) {real, imag} */,
  {32'h41ccc588, 32'hc295669b} /* (28, 16, 27) {real, imag} */,
  {32'h42ee3bee, 32'h412859de} /* (28, 16, 26) {real, imag} */,
  {32'hc20c563d, 32'hc03fe1d8} /* (28, 16, 25) {real, imag} */,
  {32'hc0d65edc, 32'hc2488308} /* (28, 16, 24) {real, imag} */,
  {32'hc1a5d242, 32'hc2ca6807} /* (28, 16, 23) {real, imag} */,
  {32'h429f2a05, 32'h41080124} /* (28, 16, 22) {real, imag} */,
  {32'h423f537d, 32'hc288d8b7} /* (28, 16, 21) {real, imag} */,
  {32'h42528722, 32'h40dd7b5e} /* (28, 16, 20) {real, imag} */,
  {32'h4277ce77, 32'hc21c89b3} /* (28, 16, 19) {real, imag} */,
  {32'hc250a208, 32'hc2870ea6} /* (28, 16, 18) {real, imag} */,
  {32'hc27186d6, 32'h4249323a} /* (28, 16, 17) {real, imag} */,
  {32'hc1c49701, 32'h00000000} /* (28, 16, 16) {real, imag} */,
  {32'hc27186d6, 32'hc249323a} /* (28, 16, 15) {real, imag} */,
  {32'hc250a208, 32'h42870ea6} /* (28, 16, 14) {real, imag} */,
  {32'h4277ce77, 32'h421c89b3} /* (28, 16, 13) {real, imag} */,
  {32'h42528722, 32'hc0dd7b5e} /* (28, 16, 12) {real, imag} */,
  {32'h423f537d, 32'h4288d8b7} /* (28, 16, 11) {real, imag} */,
  {32'h429f2a05, 32'hc1080124} /* (28, 16, 10) {real, imag} */,
  {32'hc1a5d242, 32'h42ca6807} /* (28, 16, 9) {real, imag} */,
  {32'hc0d65edc, 32'h42488308} /* (28, 16, 8) {real, imag} */,
  {32'hc20c563d, 32'h403fe1d8} /* (28, 16, 7) {real, imag} */,
  {32'h42ee3bee, 32'hc12859de} /* (28, 16, 6) {real, imag} */,
  {32'h41ccc588, 32'h4295669b} /* (28, 16, 5) {real, imag} */,
  {32'hc2a7a401, 32'hc320d283} /* (28, 16, 4) {real, imag} */,
  {32'h428e49e5, 32'hc198ffd6} /* (28, 16, 3) {real, imag} */,
  {32'h447ecd50, 32'h4345907a} /* (28, 16, 2) {real, imag} */,
  {32'hc4f21890, 32'hc3afb89e} /* (28, 16, 1) {real, imag} */,
  {32'hc4c6dd09, 32'h00000000} /* (28, 16, 0) {real, imag} */,
  {32'hc4ef3ebd, 32'h4378e370} /* (28, 15, 31) {real, imag} */,
  {32'h44837347, 32'hc37478e8} /* (28, 15, 30) {real, imag} */,
  {32'h4281cda4, 32'h41c6104b} /* (28, 15, 29) {real, imag} */,
  {32'hc3810b81, 32'h43218d38} /* (28, 15, 28) {real, imag} */,
  {32'h42ad7414, 32'hc22840ea} /* (28, 15, 27) {real, imag} */,
  {32'h42e5cf20, 32'h41c957b2} /* (28, 15, 26) {real, imag} */,
  {32'hc25d6974, 32'h41b99d05} /* (28, 15, 25) {real, imag} */,
  {32'h43126c99, 32'hc259f01e} /* (28, 15, 24) {real, imag} */,
  {32'hc1e5475c, 32'hc1b90962} /* (28, 15, 23) {real, imag} */,
  {32'hc0803110, 32'hc24d5688} /* (28, 15, 22) {real, imag} */,
  {32'h424f336f, 32'hc0294cb0} /* (28, 15, 21) {real, imag} */,
  {32'hc17d3c1a, 32'hc29f149c} /* (28, 15, 20) {real, imag} */,
  {32'hc0cfddd8, 32'hc2509315} /* (28, 15, 19) {real, imag} */,
  {32'hc17df591, 32'hc2b0bba0} /* (28, 15, 18) {real, imag} */,
  {32'h4199c662, 32'h41918268} /* (28, 15, 17) {real, imag} */,
  {32'hc23d4f56, 32'h00000000} /* (28, 15, 16) {real, imag} */,
  {32'h4199c662, 32'hc1918268} /* (28, 15, 15) {real, imag} */,
  {32'hc17df591, 32'h42b0bba0} /* (28, 15, 14) {real, imag} */,
  {32'hc0cfddd8, 32'h42509315} /* (28, 15, 13) {real, imag} */,
  {32'hc17d3c1a, 32'h429f149c} /* (28, 15, 12) {real, imag} */,
  {32'h424f336f, 32'h40294cb0} /* (28, 15, 11) {real, imag} */,
  {32'hc0803110, 32'h424d5688} /* (28, 15, 10) {real, imag} */,
  {32'hc1e5475c, 32'h41b90962} /* (28, 15, 9) {real, imag} */,
  {32'h43126c99, 32'h4259f01e} /* (28, 15, 8) {real, imag} */,
  {32'hc25d6974, 32'hc1b99d05} /* (28, 15, 7) {real, imag} */,
  {32'h42e5cf20, 32'hc1c957b2} /* (28, 15, 6) {real, imag} */,
  {32'h42ad7414, 32'h422840ea} /* (28, 15, 5) {real, imag} */,
  {32'hc3810b81, 32'hc3218d38} /* (28, 15, 4) {real, imag} */,
  {32'h4281cda4, 32'hc1c6104b} /* (28, 15, 3) {real, imag} */,
  {32'h44837347, 32'h437478e8} /* (28, 15, 2) {real, imag} */,
  {32'hc4ef3ebd, 32'hc378e370} /* (28, 15, 1) {real, imag} */,
  {32'hc4c03d80, 32'h00000000} /* (28, 15, 0) {real, imag} */,
  {32'hc4df0181, 32'h438d7108} /* (28, 14, 31) {real, imag} */,
  {32'h4478a265, 32'hc3534ee7} /* (28, 14, 30) {real, imag} */,
  {32'hc25d6a8c, 32'hc28f2214} /* (28, 14, 29) {real, imag} */,
  {32'hc3923126, 32'h4227616f} /* (28, 14, 28) {real, imag} */,
  {32'h432cd11f, 32'hc2aedc40} /* (28, 14, 27) {real, imag} */,
  {32'h4305a53f, 32'hc230f939} /* (28, 14, 26) {real, imag} */,
  {32'h41860b1d, 32'hc1c28d66} /* (28, 14, 25) {real, imag} */,
  {32'h41f1236e, 32'hc0836c90} /* (28, 14, 24) {real, imag} */,
  {32'hc2173c07, 32'hc1fbfc06} /* (28, 14, 23) {real, imag} */,
  {32'h4255b3f4, 32'hc1dc1836} /* (28, 14, 22) {real, imag} */,
  {32'hc294f967, 32'h41fc18e8} /* (28, 14, 21) {real, imag} */,
  {32'h4163bfc0, 32'hc217b84a} /* (28, 14, 20) {real, imag} */,
  {32'h41f59c1c, 32'h42055236} /* (28, 14, 19) {real, imag} */,
  {32'h4254031e, 32'hc217a7de} /* (28, 14, 18) {real, imag} */,
  {32'h4222554a, 32'hc1d93da4} /* (28, 14, 17) {real, imag} */,
  {32'h41a75a7c, 32'h00000000} /* (28, 14, 16) {real, imag} */,
  {32'h4222554a, 32'h41d93da4} /* (28, 14, 15) {real, imag} */,
  {32'h4254031e, 32'h4217a7de} /* (28, 14, 14) {real, imag} */,
  {32'h41f59c1c, 32'hc2055236} /* (28, 14, 13) {real, imag} */,
  {32'h4163bfc0, 32'h4217b84a} /* (28, 14, 12) {real, imag} */,
  {32'hc294f967, 32'hc1fc18e8} /* (28, 14, 11) {real, imag} */,
  {32'h4255b3f4, 32'h41dc1836} /* (28, 14, 10) {real, imag} */,
  {32'hc2173c07, 32'h41fbfc06} /* (28, 14, 9) {real, imag} */,
  {32'h41f1236e, 32'h40836c90} /* (28, 14, 8) {real, imag} */,
  {32'h41860b1d, 32'h41c28d66} /* (28, 14, 7) {real, imag} */,
  {32'h4305a53f, 32'h4230f939} /* (28, 14, 6) {real, imag} */,
  {32'h432cd11f, 32'h42aedc40} /* (28, 14, 5) {real, imag} */,
  {32'hc3923126, 32'hc227616f} /* (28, 14, 4) {real, imag} */,
  {32'hc25d6a8c, 32'h428f2214} /* (28, 14, 3) {real, imag} */,
  {32'h4478a265, 32'h43534ee7} /* (28, 14, 2) {real, imag} */,
  {32'hc4df0181, 32'hc38d7108} /* (28, 14, 1) {real, imag} */,
  {32'hc4ab78d7, 32'h00000000} /* (28, 14, 0) {real, imag} */,
  {32'hc4c7962a, 32'h42e8e5a2} /* (28, 13, 31) {real, imag} */,
  {32'h44443763, 32'hc1cc18e0} /* (28, 13, 30) {real, imag} */,
  {32'hc2e36ba8, 32'h419a4cb0} /* (28, 13, 29) {real, imag} */,
  {32'hc3813238, 32'hc2c1970c} /* (28, 13, 28) {real, imag} */,
  {32'h4335f20b, 32'hc2c84d8f} /* (28, 13, 27) {real, imag} */,
  {32'h429aed6b, 32'h424a7b39} /* (28, 13, 26) {real, imag} */,
  {32'h41ddb730, 32'hc1f09f90} /* (28, 13, 25) {real, imag} */,
  {32'h415c1efc, 32'hc2f55764} /* (28, 13, 24) {real, imag} */,
  {32'h4246acc8, 32'h419bef12} /* (28, 13, 23) {real, imag} */,
  {32'hc2766c08, 32'h4289ca7e} /* (28, 13, 22) {real, imag} */,
  {32'h426e5ef9, 32'h40f9858c} /* (28, 13, 21) {real, imag} */,
  {32'hc270530a, 32'hc1541578} /* (28, 13, 20) {real, imag} */,
  {32'h424e2ad7, 32'h42a85a06} /* (28, 13, 19) {real, imag} */,
  {32'hc1d90d4a, 32'h418ea850} /* (28, 13, 18) {real, imag} */,
  {32'h412c76ec, 32'hc0410090} /* (28, 13, 17) {real, imag} */,
  {32'h40f07930, 32'h00000000} /* (28, 13, 16) {real, imag} */,
  {32'h412c76ec, 32'h40410090} /* (28, 13, 15) {real, imag} */,
  {32'hc1d90d4a, 32'hc18ea850} /* (28, 13, 14) {real, imag} */,
  {32'h424e2ad7, 32'hc2a85a06} /* (28, 13, 13) {real, imag} */,
  {32'hc270530a, 32'h41541578} /* (28, 13, 12) {real, imag} */,
  {32'h426e5ef9, 32'hc0f9858c} /* (28, 13, 11) {real, imag} */,
  {32'hc2766c08, 32'hc289ca7e} /* (28, 13, 10) {real, imag} */,
  {32'h4246acc8, 32'hc19bef12} /* (28, 13, 9) {real, imag} */,
  {32'h415c1efc, 32'h42f55764} /* (28, 13, 8) {real, imag} */,
  {32'h41ddb730, 32'h41f09f90} /* (28, 13, 7) {real, imag} */,
  {32'h429aed6b, 32'hc24a7b39} /* (28, 13, 6) {real, imag} */,
  {32'h4335f20b, 32'h42c84d8f} /* (28, 13, 5) {real, imag} */,
  {32'hc3813238, 32'h42c1970c} /* (28, 13, 4) {real, imag} */,
  {32'hc2e36ba8, 32'hc19a4cb0} /* (28, 13, 3) {real, imag} */,
  {32'h44443763, 32'h41cc18e0} /* (28, 13, 2) {real, imag} */,
  {32'hc4c7962a, 32'hc2e8e5a2} /* (28, 13, 1) {real, imag} */,
  {32'hc4976e22, 32'h00000000} /* (28, 13, 0) {real, imag} */,
  {32'hc4b4db04, 32'h4307d650} /* (28, 12, 31) {real, imag} */,
  {32'h4413bc86, 32'hc115d170} /* (28, 12, 30) {real, imag} */,
  {32'hbe8cf200, 32'hc3030e43} /* (28, 12, 29) {real, imag} */,
  {32'hc30c745a, 32'hc2678978} /* (28, 12, 28) {real, imag} */,
  {32'h43238b1c, 32'hc335dbff} /* (28, 12, 27) {real, imag} */,
  {32'h41a691c9, 32'h41210eb6} /* (28, 12, 26) {real, imag} */,
  {32'h4291d1d4, 32'h42090661} /* (28, 12, 25) {real, imag} */,
  {32'h428cb1a6, 32'hc2982250} /* (28, 12, 24) {real, imag} */,
  {32'h41db282c, 32'hc2c2c39c} /* (28, 12, 23) {real, imag} */,
  {32'hc1c43e18, 32'hc23ce560} /* (28, 12, 22) {real, imag} */,
  {32'hc0863060, 32'hc2a69c13} /* (28, 12, 21) {real, imag} */,
  {32'hc19a43ce, 32'hc24d4afa} /* (28, 12, 20) {real, imag} */,
  {32'h416f1664, 32'hc2559726} /* (28, 12, 19) {real, imag} */,
  {32'h424657ec, 32'hc2f82a74} /* (28, 12, 18) {real, imag} */,
  {32'hc21a1615, 32'hc1be6ab4} /* (28, 12, 17) {real, imag} */,
  {32'h419f3d67, 32'h00000000} /* (28, 12, 16) {real, imag} */,
  {32'hc21a1615, 32'h41be6ab4} /* (28, 12, 15) {real, imag} */,
  {32'h424657ec, 32'h42f82a74} /* (28, 12, 14) {real, imag} */,
  {32'h416f1664, 32'h42559726} /* (28, 12, 13) {real, imag} */,
  {32'hc19a43ce, 32'h424d4afa} /* (28, 12, 12) {real, imag} */,
  {32'hc0863060, 32'h42a69c13} /* (28, 12, 11) {real, imag} */,
  {32'hc1c43e18, 32'h423ce560} /* (28, 12, 10) {real, imag} */,
  {32'h41db282c, 32'h42c2c39c} /* (28, 12, 9) {real, imag} */,
  {32'h428cb1a6, 32'h42982250} /* (28, 12, 8) {real, imag} */,
  {32'h4291d1d4, 32'hc2090661} /* (28, 12, 7) {real, imag} */,
  {32'h41a691c9, 32'hc1210eb6} /* (28, 12, 6) {real, imag} */,
  {32'h43238b1c, 32'h4335dbff} /* (28, 12, 5) {real, imag} */,
  {32'hc30c745a, 32'h42678978} /* (28, 12, 4) {real, imag} */,
  {32'hbe8cf200, 32'h43030e43} /* (28, 12, 3) {real, imag} */,
  {32'h4413bc86, 32'h4115d170} /* (28, 12, 2) {real, imag} */,
  {32'hc4b4db04, 32'hc307d650} /* (28, 12, 1) {real, imag} */,
  {32'hc49b57a8, 32'h00000000} /* (28, 12, 0) {real, imag} */,
  {32'hc43eb820, 32'h42a06d2a} /* (28, 11, 31) {real, imag} */,
  {32'h43de82ce, 32'hc28345b0} /* (28, 11, 30) {real, imag} */,
  {32'h40dc3b9c, 32'hc227308e} /* (28, 11, 29) {real, imag} */,
  {32'hc2859845, 32'hc278c801} /* (28, 11, 28) {real, imag} */,
  {32'h41953f4e, 32'hc284e476} /* (28, 11, 27) {real, imag} */,
  {32'hc2befd8a, 32'hc250cd42} /* (28, 11, 26) {real, imag} */,
  {32'h4194b5a8, 32'hc2be9d58} /* (28, 11, 25) {real, imag} */,
  {32'h42ac4636, 32'h4243bbc2} /* (28, 11, 24) {real, imag} */,
  {32'h427b2c22, 32'h42323078} /* (28, 11, 23) {real, imag} */,
  {32'h4274339b, 32'h41c5f6f2} /* (28, 11, 22) {real, imag} */,
  {32'h4138b741, 32'hc11677b0} /* (28, 11, 21) {real, imag} */,
  {32'h4114fbd4, 32'h42967ecb} /* (28, 11, 20) {real, imag} */,
  {32'hc274e0d8, 32'h40bc5ee0} /* (28, 11, 19) {real, imag} */,
  {32'hc075fd30, 32'hc0377bc0} /* (28, 11, 18) {real, imag} */,
  {32'h42206d99, 32'hc034d078} /* (28, 11, 17) {real, imag} */,
  {32'hc2c9a405, 32'h00000000} /* (28, 11, 16) {real, imag} */,
  {32'h42206d99, 32'h4034d078} /* (28, 11, 15) {real, imag} */,
  {32'hc075fd30, 32'h40377bc0} /* (28, 11, 14) {real, imag} */,
  {32'hc274e0d8, 32'hc0bc5ee0} /* (28, 11, 13) {real, imag} */,
  {32'h4114fbd4, 32'hc2967ecb} /* (28, 11, 12) {real, imag} */,
  {32'h4138b741, 32'h411677b0} /* (28, 11, 11) {real, imag} */,
  {32'h4274339b, 32'hc1c5f6f2} /* (28, 11, 10) {real, imag} */,
  {32'h427b2c22, 32'hc2323078} /* (28, 11, 9) {real, imag} */,
  {32'h42ac4636, 32'hc243bbc2} /* (28, 11, 8) {real, imag} */,
  {32'h4194b5a8, 32'h42be9d58} /* (28, 11, 7) {real, imag} */,
  {32'hc2befd8a, 32'h4250cd42} /* (28, 11, 6) {real, imag} */,
  {32'h41953f4e, 32'h4284e476} /* (28, 11, 5) {real, imag} */,
  {32'hc2859845, 32'h4278c801} /* (28, 11, 4) {real, imag} */,
  {32'h40dc3b9c, 32'h4227308e} /* (28, 11, 3) {real, imag} */,
  {32'h43de82ce, 32'h428345b0} /* (28, 11, 2) {real, imag} */,
  {32'hc43eb820, 32'hc2a06d2a} /* (28, 11, 1) {real, imag} */,
  {32'hc460886c, 32'h00000000} /* (28, 11, 0) {real, imag} */,
  {32'h43c9b7dc, 32'hc2c91ca1} /* (28, 10, 31) {real, imag} */,
  {32'hc38e77e4, 32'h42d50bd2} /* (28, 10, 30) {real, imag} */,
  {32'h41b43350, 32'h42c110b9} /* (28, 10, 29) {real, imag} */,
  {32'h4353203c, 32'hc33a4392} /* (28, 10, 28) {real, imag} */,
  {32'hc30103f2, 32'hc20778b1} /* (28, 10, 27) {real, imag} */,
  {32'hc1e6e4e5, 32'hc0fecd7c} /* (28, 10, 26) {real, imag} */,
  {32'h42df19ec, 32'hbfabac00} /* (28, 10, 25) {real, imag} */,
  {32'hc19af524, 32'h41d5491e} /* (28, 10, 24) {real, imag} */,
  {32'hc1c57af5, 32'h416f731c} /* (28, 10, 23) {real, imag} */,
  {32'hc09d405c, 32'hc2c4e615} /* (28, 10, 22) {real, imag} */,
  {32'hc300e845, 32'h429ebc12} /* (28, 10, 21) {real, imag} */,
  {32'h42cbc56b, 32'hc24b2c8c} /* (28, 10, 20) {real, imag} */,
  {32'h40962994, 32'h416168c0} /* (28, 10, 19) {real, imag} */,
  {32'hc1c59203, 32'hc10b75a0} /* (28, 10, 18) {real, imag} */,
  {32'h40836adc, 32'h422409a5} /* (28, 10, 17) {real, imag} */,
  {32'hc101f1bc, 32'h00000000} /* (28, 10, 16) {real, imag} */,
  {32'h40836adc, 32'hc22409a5} /* (28, 10, 15) {real, imag} */,
  {32'hc1c59203, 32'h410b75a0} /* (28, 10, 14) {real, imag} */,
  {32'h40962994, 32'hc16168c0} /* (28, 10, 13) {real, imag} */,
  {32'h42cbc56b, 32'h424b2c8c} /* (28, 10, 12) {real, imag} */,
  {32'hc300e845, 32'hc29ebc12} /* (28, 10, 11) {real, imag} */,
  {32'hc09d405c, 32'h42c4e615} /* (28, 10, 10) {real, imag} */,
  {32'hc1c57af5, 32'hc16f731c} /* (28, 10, 9) {real, imag} */,
  {32'hc19af524, 32'hc1d5491e} /* (28, 10, 8) {real, imag} */,
  {32'h42df19ec, 32'h3fabac00} /* (28, 10, 7) {real, imag} */,
  {32'hc1e6e4e5, 32'h40fecd7c} /* (28, 10, 6) {real, imag} */,
  {32'hc30103f2, 32'h420778b1} /* (28, 10, 5) {real, imag} */,
  {32'h4353203c, 32'h433a4392} /* (28, 10, 4) {real, imag} */,
  {32'h41b43350, 32'hc2c110b9} /* (28, 10, 3) {real, imag} */,
  {32'hc38e77e4, 32'hc2d50bd2} /* (28, 10, 2) {real, imag} */,
  {32'h43c9b7dc, 32'h42c91ca1} /* (28, 10, 1) {real, imag} */,
  {32'hc29e9ec8, 32'h00000000} /* (28, 10, 0) {real, imag} */,
  {32'h448feaa6, 32'hc2fa4f92} /* (28, 9, 31) {real, imag} */,
  {32'hc41fa5be, 32'h4317a9df} /* (28, 9, 30) {real, imag} */,
  {32'h42fa53d0, 32'h42d17d4f} /* (28, 9, 29) {real, imag} */,
  {32'h4317f8d5, 32'hc3327a1c} /* (28, 9, 28) {real, imag} */,
  {32'hc3569f8d, 32'h424a829c} /* (28, 9, 27) {real, imag} */,
  {32'hc2bdbd44, 32'hc31e8720} /* (28, 9, 26) {real, imag} */,
  {32'h42b0eb49, 32'hc2652418} /* (28, 9, 25) {real, imag} */,
  {32'hc290c9f6, 32'h41ee3b08} /* (28, 9, 24) {real, imag} */,
  {32'h4235a4e1, 32'hc227a0f8} /* (28, 9, 23) {real, imag} */,
  {32'hbfd43cc0, 32'hc2db7d56} /* (28, 9, 22) {real, imag} */,
  {32'hc2b3ae2f, 32'h431cc365} /* (28, 9, 21) {real, imag} */,
  {32'h40f28e20, 32'hc0ce06fc} /* (28, 9, 20) {real, imag} */,
  {32'hc1dcb383, 32'hc1677d4c} /* (28, 9, 19) {real, imag} */,
  {32'h41dba9fe, 32'hc24fc501} /* (28, 9, 18) {real, imag} */,
  {32'hc1ed7876, 32'hc112ac04} /* (28, 9, 17) {real, imag} */,
  {32'hc1c8e472, 32'h00000000} /* (28, 9, 16) {real, imag} */,
  {32'hc1ed7876, 32'h4112ac04} /* (28, 9, 15) {real, imag} */,
  {32'h41dba9fe, 32'h424fc501} /* (28, 9, 14) {real, imag} */,
  {32'hc1dcb383, 32'h41677d4c} /* (28, 9, 13) {real, imag} */,
  {32'h40f28e20, 32'h40ce06fc} /* (28, 9, 12) {real, imag} */,
  {32'hc2b3ae2f, 32'hc31cc365} /* (28, 9, 11) {real, imag} */,
  {32'hbfd43cc0, 32'h42db7d56} /* (28, 9, 10) {real, imag} */,
  {32'h4235a4e1, 32'h4227a0f8} /* (28, 9, 9) {real, imag} */,
  {32'hc290c9f6, 32'hc1ee3b08} /* (28, 9, 8) {real, imag} */,
  {32'h42b0eb49, 32'h42652418} /* (28, 9, 7) {real, imag} */,
  {32'hc2bdbd44, 32'h431e8720} /* (28, 9, 6) {real, imag} */,
  {32'hc3569f8d, 32'hc24a829c} /* (28, 9, 5) {real, imag} */,
  {32'h4317f8d5, 32'h43327a1c} /* (28, 9, 4) {real, imag} */,
  {32'h42fa53d0, 32'hc2d17d4f} /* (28, 9, 3) {real, imag} */,
  {32'hc41fa5be, 32'hc317a9df} /* (28, 9, 2) {real, imag} */,
  {32'h448feaa6, 32'h42fa4f92} /* (28, 9, 1) {real, imag} */,
  {32'h43ffed35, 32'h00000000} /* (28, 9, 0) {real, imag} */,
  {32'h44b1c2b4, 32'hc338f064} /* (28, 8, 31) {real, imag} */,
  {32'hc41b3104, 32'h4393a8ea} /* (28, 8, 30) {real, imag} */,
  {32'h43169538, 32'h425f7da0} /* (28, 8, 29) {real, imag} */,
  {32'h43209392, 32'hc2a8e2c8} /* (28, 8, 28) {real, imag} */,
  {32'hc31a6813, 32'h4339165b} /* (28, 8, 27) {real, imag} */,
  {32'h425051ac, 32'hc2cc033c} /* (28, 8, 26) {real, imag} */,
  {32'hc2446596, 32'h41f97458} /* (28, 8, 25) {real, imag} */,
  {32'hc265bf04, 32'h418d3fd4} /* (28, 8, 24) {real, imag} */,
  {32'hc2b480d1, 32'h424e49fa} /* (28, 8, 23) {real, imag} */,
  {32'h42e7094a, 32'hc0ab2cae} /* (28, 8, 22) {real, imag} */,
  {32'hbfa21e80, 32'h42103fa4} /* (28, 8, 21) {real, imag} */,
  {32'hc237f355, 32'hc25f984b} /* (28, 8, 20) {real, imag} */,
  {32'h418a59b0, 32'hc2bcfc58} /* (28, 8, 19) {real, imag} */,
  {32'hc2b792a2, 32'h42712bd2} /* (28, 8, 18) {real, imag} */,
  {32'hc1f0c014, 32'h404bfc10} /* (28, 8, 17) {real, imag} */,
  {32'hc1e35c03, 32'h00000000} /* (28, 8, 16) {real, imag} */,
  {32'hc1f0c014, 32'hc04bfc10} /* (28, 8, 15) {real, imag} */,
  {32'hc2b792a2, 32'hc2712bd2} /* (28, 8, 14) {real, imag} */,
  {32'h418a59b0, 32'h42bcfc58} /* (28, 8, 13) {real, imag} */,
  {32'hc237f355, 32'h425f984b} /* (28, 8, 12) {real, imag} */,
  {32'hbfa21e80, 32'hc2103fa4} /* (28, 8, 11) {real, imag} */,
  {32'h42e7094a, 32'h40ab2cae} /* (28, 8, 10) {real, imag} */,
  {32'hc2b480d1, 32'hc24e49fa} /* (28, 8, 9) {real, imag} */,
  {32'hc265bf04, 32'hc18d3fd4} /* (28, 8, 8) {real, imag} */,
  {32'hc2446596, 32'hc1f97458} /* (28, 8, 7) {real, imag} */,
  {32'h425051ac, 32'h42cc033c} /* (28, 8, 6) {real, imag} */,
  {32'hc31a6813, 32'hc339165b} /* (28, 8, 5) {real, imag} */,
  {32'h43209392, 32'h42a8e2c8} /* (28, 8, 4) {real, imag} */,
  {32'h43169538, 32'hc25f7da0} /* (28, 8, 3) {real, imag} */,
  {32'hc41b3104, 32'hc393a8ea} /* (28, 8, 2) {real, imag} */,
  {32'h44b1c2b4, 32'h4338f064} /* (28, 8, 1) {real, imag} */,
  {32'h43f993e8, 32'h00000000} /* (28, 8, 0) {real, imag} */,
  {32'h44ba4d48, 32'hc379e26d} /* (28, 7, 31) {real, imag} */,
  {32'hc4308cc3, 32'h43d5dc22} /* (28, 7, 30) {real, imag} */,
  {32'h40ff50f0, 32'h433c75ce} /* (28, 7, 29) {real, imag} */,
  {32'h4321db47, 32'hc205613c} /* (28, 7, 28) {real, imag} */,
  {32'hc3144ffb, 32'h40ee7e80} /* (28, 7, 27) {real, imag} */,
  {32'hc26fcee1, 32'hc2051b5e} /* (28, 7, 26) {real, imag} */,
  {32'hc273d22d, 32'hc2a9c3a0} /* (28, 7, 25) {real, imag} */,
  {32'hc14b3cf2, 32'h42d3890e} /* (28, 7, 24) {real, imag} */,
  {32'h418a9286, 32'hbf3bd580} /* (28, 7, 23) {real, imag} */,
  {32'hc2f80265, 32'hc131a52c} /* (28, 7, 22) {real, imag} */,
  {32'hc249cd06, 32'h426e98df} /* (28, 7, 21) {real, imag} */,
  {32'h42ec69a6, 32'hc2429722} /* (28, 7, 20) {real, imag} */,
  {32'hc2996740, 32'hc171788c} /* (28, 7, 19) {real, imag} */,
  {32'h4283c608, 32'h411b606e} /* (28, 7, 18) {real, imag} */,
  {32'hc25c313a, 32'h41cbe8ee} /* (28, 7, 17) {real, imag} */,
  {32'h42ad69be, 32'h00000000} /* (28, 7, 16) {real, imag} */,
  {32'hc25c313a, 32'hc1cbe8ee} /* (28, 7, 15) {real, imag} */,
  {32'h4283c608, 32'hc11b606e} /* (28, 7, 14) {real, imag} */,
  {32'hc2996740, 32'h4171788c} /* (28, 7, 13) {real, imag} */,
  {32'h42ec69a6, 32'h42429722} /* (28, 7, 12) {real, imag} */,
  {32'hc249cd06, 32'hc26e98df} /* (28, 7, 11) {real, imag} */,
  {32'hc2f80265, 32'h4131a52c} /* (28, 7, 10) {real, imag} */,
  {32'h418a9286, 32'h3f3bd580} /* (28, 7, 9) {real, imag} */,
  {32'hc14b3cf2, 32'hc2d3890e} /* (28, 7, 8) {real, imag} */,
  {32'hc273d22d, 32'h42a9c3a0} /* (28, 7, 7) {real, imag} */,
  {32'hc26fcee1, 32'h42051b5e} /* (28, 7, 6) {real, imag} */,
  {32'hc3144ffb, 32'hc0ee7e80} /* (28, 7, 5) {real, imag} */,
  {32'h4321db47, 32'h4205613c} /* (28, 7, 4) {real, imag} */,
  {32'h40ff50f0, 32'hc33c75ce} /* (28, 7, 3) {real, imag} */,
  {32'hc4308cc3, 32'hc3d5dc22} /* (28, 7, 2) {real, imag} */,
  {32'h44ba4d48, 32'h4379e26d} /* (28, 7, 1) {real, imag} */,
  {32'h43fc9073, 32'h00000000} /* (28, 7, 0) {real, imag} */,
  {32'h44a9b921, 32'hc3dc5ba1} /* (28, 6, 31) {real, imag} */,
  {32'hc4244ea2, 32'h4409926d} /* (28, 6, 30) {real, imag} */,
  {32'hc2b670a6, 32'h42cd7419} /* (28, 6, 29) {real, imag} */,
  {32'h40787160, 32'hc08e0410} /* (28, 6, 28) {real, imag} */,
  {32'hc37ab7bf, 32'h41e41880} /* (28, 6, 27) {real, imag} */,
  {32'h42d85c96, 32'hc30964ee} /* (28, 6, 26) {real, imag} */,
  {32'hc08a5bb8, 32'hc32e30f4} /* (28, 6, 25) {real, imag} */,
  {32'hc103c025, 32'h422a498a} /* (28, 6, 24) {real, imag} */,
  {32'h42aea39f, 32'h42649ddf} /* (28, 6, 23) {real, imag} */,
  {32'h4244c35e, 32'h420ad18e} /* (28, 6, 22) {real, imag} */,
  {32'hc20a4d7c, 32'hc0981d9c} /* (28, 6, 21) {real, imag} */,
  {32'hc24aaffe, 32'hc00d85f8} /* (28, 6, 20) {real, imag} */,
  {32'hc2034170, 32'hc1b78c2e} /* (28, 6, 19) {real, imag} */,
  {32'hc1990f98, 32'hc259d0e7} /* (28, 6, 18) {real, imag} */,
  {32'h413bc7c0, 32'hc2163804} /* (28, 6, 17) {real, imag} */,
  {32'hc0a48c44, 32'h00000000} /* (28, 6, 16) {real, imag} */,
  {32'h413bc7c0, 32'h42163804} /* (28, 6, 15) {real, imag} */,
  {32'hc1990f98, 32'h4259d0e7} /* (28, 6, 14) {real, imag} */,
  {32'hc2034170, 32'h41b78c2e} /* (28, 6, 13) {real, imag} */,
  {32'hc24aaffe, 32'h400d85f8} /* (28, 6, 12) {real, imag} */,
  {32'hc20a4d7c, 32'h40981d9c} /* (28, 6, 11) {real, imag} */,
  {32'h4244c35e, 32'hc20ad18e} /* (28, 6, 10) {real, imag} */,
  {32'h42aea39f, 32'hc2649ddf} /* (28, 6, 9) {real, imag} */,
  {32'hc103c025, 32'hc22a498a} /* (28, 6, 8) {real, imag} */,
  {32'hc08a5bb8, 32'h432e30f4} /* (28, 6, 7) {real, imag} */,
  {32'h42d85c96, 32'h430964ee} /* (28, 6, 6) {real, imag} */,
  {32'hc37ab7bf, 32'hc1e41880} /* (28, 6, 5) {real, imag} */,
  {32'h40787160, 32'h408e0410} /* (28, 6, 4) {real, imag} */,
  {32'hc2b670a6, 32'hc2cd7419} /* (28, 6, 3) {real, imag} */,
  {32'hc4244ea2, 32'hc409926d} /* (28, 6, 2) {real, imag} */,
  {32'h44a9b921, 32'h43dc5ba1} /* (28, 6, 1) {real, imag} */,
  {32'h441b7c22, 32'h00000000} /* (28, 6, 0) {real, imag} */,
  {32'h4472f530, 32'hc46f78f7} /* (28, 5, 31) {real, imag} */,
  {32'hc3745edc, 32'h443a0623} /* (28, 5, 30) {real, imag} */,
  {32'hc3002d79, 32'h422ff21e} /* (28, 5, 29) {real, imag} */,
  {32'hc2a00f74, 32'h4207d995} /* (28, 5, 28) {real, imag} */,
  {32'hc2f7e18a, 32'h42327eba} /* (28, 5, 27) {real, imag} */,
  {32'h41676aac, 32'hc2cb9469} /* (28, 5, 26) {real, imag} */,
  {32'h41abb09a, 32'hc221de39} /* (28, 5, 25) {real, imag} */,
  {32'h42a823f3, 32'h4252293e} /* (28, 5, 24) {real, imag} */,
  {32'hc266b57e, 32'h421e7c71} /* (28, 5, 23) {real, imag} */,
  {32'hc2a093b2, 32'hc221ad58} /* (28, 5, 22) {real, imag} */,
  {32'h42b4aade, 32'h4239f914} /* (28, 5, 21) {real, imag} */,
  {32'h3fe2b5dc, 32'hc1c0e5f8} /* (28, 5, 20) {real, imag} */,
  {32'h424278c6, 32'h40eb7940} /* (28, 5, 19) {real, imag} */,
  {32'h41923a08, 32'h4280bb48} /* (28, 5, 18) {real, imag} */,
  {32'hc2212d4a, 32'hc12b2448} /* (28, 5, 17) {real, imag} */,
  {32'hc2108a04, 32'h00000000} /* (28, 5, 16) {real, imag} */,
  {32'hc2212d4a, 32'h412b2448} /* (28, 5, 15) {real, imag} */,
  {32'h41923a08, 32'hc280bb48} /* (28, 5, 14) {real, imag} */,
  {32'h424278c6, 32'hc0eb7940} /* (28, 5, 13) {real, imag} */,
  {32'h3fe2b5dc, 32'h41c0e5f8} /* (28, 5, 12) {real, imag} */,
  {32'h42b4aade, 32'hc239f914} /* (28, 5, 11) {real, imag} */,
  {32'hc2a093b2, 32'h4221ad58} /* (28, 5, 10) {real, imag} */,
  {32'hc266b57e, 32'hc21e7c71} /* (28, 5, 9) {real, imag} */,
  {32'h42a823f3, 32'hc252293e} /* (28, 5, 8) {real, imag} */,
  {32'h41abb09a, 32'h4221de39} /* (28, 5, 7) {real, imag} */,
  {32'h41676aac, 32'h42cb9469} /* (28, 5, 6) {real, imag} */,
  {32'hc2f7e18a, 32'hc2327eba} /* (28, 5, 5) {real, imag} */,
  {32'hc2a00f74, 32'hc207d995} /* (28, 5, 4) {real, imag} */,
  {32'hc3002d79, 32'hc22ff21e} /* (28, 5, 3) {real, imag} */,
  {32'hc3745edc, 32'hc43a0623} /* (28, 5, 2) {real, imag} */,
  {32'h4472f530, 32'h446f78f7} /* (28, 5, 1) {real, imag} */,
  {32'h44371df0, 32'h00000000} /* (28, 5, 0) {real, imag} */,
  {32'h441481cf, 32'hc47dd97e} /* (28, 4, 31) {real, imag} */,
  {32'h43731362, 32'h44417651} /* (28, 4, 30) {real, imag} */,
  {32'hc292c620, 32'hc2850a8b} /* (28, 4, 29) {real, imag} */,
  {32'hc30dce06, 32'h42bfb086} /* (28, 4, 28) {real, imag} */,
  {32'hc3802238, 32'hc2c097e2} /* (28, 4, 27) {real, imag} */,
  {32'hc29e7926, 32'h42c6a92d} /* (28, 4, 26) {real, imag} */,
  {32'h41b5559c, 32'hc273288a} /* (28, 4, 25) {real, imag} */,
  {32'h4241908f, 32'h42442de5} /* (28, 4, 24) {real, imag} */,
  {32'hc2804763, 32'hc20f2a1a} /* (28, 4, 23) {real, imag} */,
  {32'hc2d50bfa, 32'hc1e8352c} /* (28, 4, 22) {real, imag} */,
  {32'h41b4989c, 32'h417961b8} /* (28, 4, 21) {real, imag} */,
  {32'h4213a655, 32'hc20c23a7} /* (28, 4, 20) {real, imag} */,
  {32'hc1c2322d, 32'hc2d7d7e3} /* (28, 4, 19) {real, imag} */,
  {32'h42855b2d, 32'h424924b0} /* (28, 4, 18) {real, imag} */,
  {32'h3eb82580, 32'h41077248} /* (28, 4, 17) {real, imag} */,
  {32'h40e1be68, 32'h00000000} /* (28, 4, 16) {real, imag} */,
  {32'h3eb82580, 32'hc1077248} /* (28, 4, 15) {real, imag} */,
  {32'h42855b2d, 32'hc24924b0} /* (28, 4, 14) {real, imag} */,
  {32'hc1c2322d, 32'h42d7d7e3} /* (28, 4, 13) {real, imag} */,
  {32'h4213a655, 32'h420c23a7} /* (28, 4, 12) {real, imag} */,
  {32'h41b4989c, 32'hc17961b8} /* (28, 4, 11) {real, imag} */,
  {32'hc2d50bfa, 32'h41e8352c} /* (28, 4, 10) {real, imag} */,
  {32'hc2804763, 32'h420f2a1a} /* (28, 4, 9) {real, imag} */,
  {32'h4241908f, 32'hc2442de5} /* (28, 4, 8) {real, imag} */,
  {32'h41b5559c, 32'h4273288a} /* (28, 4, 7) {real, imag} */,
  {32'hc29e7926, 32'hc2c6a92d} /* (28, 4, 6) {real, imag} */,
  {32'hc3802238, 32'h42c097e2} /* (28, 4, 5) {real, imag} */,
  {32'hc30dce06, 32'hc2bfb086} /* (28, 4, 4) {real, imag} */,
  {32'hc292c620, 32'h42850a8b} /* (28, 4, 3) {real, imag} */,
  {32'h43731362, 32'hc4417651} /* (28, 4, 2) {real, imag} */,
  {32'h441481cf, 32'h447dd97e} /* (28, 4, 1) {real, imag} */,
  {32'h43eab082, 32'h00000000} /* (28, 4, 0) {real, imag} */,
  {32'h43fc6528, 32'hc49529fc} /* (28, 3, 31) {real, imag} */,
  {32'h43d6ad28, 32'h4423b55e} /* (28, 3, 30) {real, imag} */,
  {32'hc2e4beb7, 32'hc30a5510} /* (28, 3, 29) {real, imag} */,
  {32'hc2f7fd9b, 32'h438bfef8} /* (28, 3, 28) {real, imag} */,
  {32'hc3808ee1, 32'h42e1232d} /* (28, 3, 27) {real, imag} */,
  {32'hc10f86fe, 32'h431a0b38} /* (28, 3, 26) {real, imag} */,
  {32'hc2a9012e, 32'hc240ec12} /* (28, 3, 25) {real, imag} */,
  {32'h420cbdda, 32'hc2462967} /* (28, 3, 24) {real, imag} */,
  {32'hc181e1a4, 32'hc22f88f6} /* (28, 3, 23) {real, imag} */,
  {32'hc188d4dc, 32'h428f131f} /* (28, 3, 22) {real, imag} */,
  {32'hc2a10e24, 32'hc2921858} /* (28, 3, 21) {real, imag} */,
  {32'hc1cec0e2, 32'hc187b56a} /* (28, 3, 20) {real, imag} */,
  {32'hc18f1b73, 32'h40d32c68} /* (28, 3, 19) {real, imag} */,
  {32'h429157d6, 32'hc18a4fd9} /* (28, 3, 18) {real, imag} */,
  {32'hc165541b, 32'h426548ce} /* (28, 3, 17) {real, imag} */,
  {32'h4180b9ee, 32'h00000000} /* (28, 3, 16) {real, imag} */,
  {32'hc165541b, 32'hc26548ce} /* (28, 3, 15) {real, imag} */,
  {32'h429157d6, 32'h418a4fd9} /* (28, 3, 14) {real, imag} */,
  {32'hc18f1b73, 32'hc0d32c68} /* (28, 3, 13) {real, imag} */,
  {32'hc1cec0e2, 32'h4187b56a} /* (28, 3, 12) {real, imag} */,
  {32'hc2a10e24, 32'h42921858} /* (28, 3, 11) {real, imag} */,
  {32'hc188d4dc, 32'hc28f131f} /* (28, 3, 10) {real, imag} */,
  {32'hc181e1a4, 32'h422f88f6} /* (28, 3, 9) {real, imag} */,
  {32'h420cbdda, 32'h42462967} /* (28, 3, 8) {real, imag} */,
  {32'hc2a9012e, 32'h4240ec12} /* (28, 3, 7) {real, imag} */,
  {32'hc10f86fe, 32'hc31a0b38} /* (28, 3, 6) {real, imag} */,
  {32'hc3808ee1, 32'hc2e1232d} /* (28, 3, 5) {real, imag} */,
  {32'hc2f7fd9b, 32'hc38bfef8} /* (28, 3, 4) {real, imag} */,
  {32'hc2e4beb7, 32'h430a5510} /* (28, 3, 3) {real, imag} */,
  {32'h43d6ad28, 32'hc423b55e} /* (28, 3, 2) {real, imag} */,
  {32'h43fc6528, 32'h449529fc} /* (28, 3, 1) {real, imag} */,
  {32'h43ee52b9, 32'h00000000} /* (28, 3, 0) {real, imag} */,
  {32'h43e045eb, 32'hc4b33540} /* (28, 2, 31) {real, imag} */,
  {32'h43a24e4e, 32'h443a4f90} /* (28, 2, 30) {real, imag} */,
  {32'hc1a1c890, 32'h42690570} /* (28, 2, 29) {real, imag} */,
  {32'hc2f8d4fe, 32'h430aa7ce} /* (28, 2, 28) {real, imag} */,
  {32'hc263d697, 32'hc2809f84} /* (28, 2, 27) {real, imag} */,
  {32'hc1f59fc8, 32'h42e7c2ec} /* (28, 2, 26) {real, imag} */,
  {32'hc341f8a0, 32'hc1ea8efa} /* (28, 2, 25) {real, imag} */,
  {32'h43135e58, 32'hc2f49e50} /* (28, 2, 24) {real, imag} */,
  {32'hc22fc5b4, 32'h40a7d866} /* (28, 2, 23) {real, imag} */,
  {32'hc20de586, 32'h430a3439} /* (28, 2, 22) {real, imag} */,
  {32'hc1df5364, 32'hc22e98fe} /* (28, 2, 21) {real, imag} */,
  {32'h42d28704, 32'h42b5bed4} /* (28, 2, 20) {real, imag} */,
  {32'h4184bd5e, 32'h41abaf96} /* (28, 2, 19) {real, imag} */,
  {32'h4133ac32, 32'h3fa131b0} /* (28, 2, 18) {real, imag} */,
  {32'hc27c7400, 32'h4201cba2} /* (28, 2, 17) {real, imag} */,
  {32'h429cf039, 32'h00000000} /* (28, 2, 16) {real, imag} */,
  {32'hc27c7400, 32'hc201cba2} /* (28, 2, 15) {real, imag} */,
  {32'h4133ac32, 32'hbfa131b0} /* (28, 2, 14) {real, imag} */,
  {32'h4184bd5e, 32'hc1abaf96} /* (28, 2, 13) {real, imag} */,
  {32'h42d28704, 32'hc2b5bed4} /* (28, 2, 12) {real, imag} */,
  {32'hc1df5364, 32'h422e98fe} /* (28, 2, 11) {real, imag} */,
  {32'hc20de586, 32'hc30a3439} /* (28, 2, 10) {real, imag} */,
  {32'hc22fc5b4, 32'hc0a7d866} /* (28, 2, 9) {real, imag} */,
  {32'h43135e58, 32'h42f49e50} /* (28, 2, 8) {real, imag} */,
  {32'hc341f8a0, 32'h41ea8efa} /* (28, 2, 7) {real, imag} */,
  {32'hc1f59fc8, 32'hc2e7c2ec} /* (28, 2, 6) {real, imag} */,
  {32'hc263d697, 32'h42809f84} /* (28, 2, 5) {real, imag} */,
  {32'hc2f8d4fe, 32'hc30aa7ce} /* (28, 2, 4) {real, imag} */,
  {32'hc1a1c890, 32'hc2690570} /* (28, 2, 3) {real, imag} */,
  {32'h43a24e4e, 32'hc43a4f90} /* (28, 2, 2) {real, imag} */,
  {32'h43e045eb, 32'h44b33540} /* (28, 2, 1) {real, imag} */,
  {32'h437ff914, 32'h00000000} /* (28, 2, 0) {real, imag} */,
  {32'h437c1e36, 32'hc4a45798} /* (28, 1, 31) {real, imag} */,
  {32'h438e691d, 32'h445a6975} /* (28, 1, 30) {real, imag} */,
  {32'hc29ca86c, 32'h41666372} /* (28, 1, 29) {real, imag} */,
  {32'h41fcee46, 32'h429caf3e} /* (28, 1, 28) {real, imag} */,
  {32'hc3539d83, 32'hc2f76442} /* (28, 1, 27) {real, imag} */,
  {32'hc10ba4d6, 32'h4332fd9c} /* (28, 1, 26) {real, imag} */,
  {32'hc2676a1b, 32'hc2b09d02} /* (28, 1, 25) {real, imag} */,
  {32'h41f20306, 32'hc29e6c5a} /* (28, 1, 24) {real, imag} */,
  {32'h4223836c, 32'h42669cff} /* (28, 1, 23) {real, imag} */,
  {32'hc2b2b54e, 32'h426197d0} /* (28, 1, 22) {real, imag} */,
  {32'h41974e47, 32'hc2849da7} /* (28, 1, 21) {real, imag} */,
  {32'h42e2ac7b, 32'h41140054} /* (28, 1, 20) {real, imag} */,
  {32'hc2ca8720, 32'hc194a3bf} /* (28, 1, 19) {real, imag} */,
  {32'h3fd92060, 32'hc1a27e02} /* (28, 1, 18) {real, imag} */,
  {32'hc202228e, 32'hc278762a} /* (28, 1, 17) {real, imag} */,
  {32'hc1041756, 32'h00000000} /* (28, 1, 16) {real, imag} */,
  {32'hc202228e, 32'h4278762a} /* (28, 1, 15) {real, imag} */,
  {32'h3fd92060, 32'h41a27e02} /* (28, 1, 14) {real, imag} */,
  {32'hc2ca8720, 32'h4194a3bf} /* (28, 1, 13) {real, imag} */,
  {32'h42e2ac7b, 32'hc1140054} /* (28, 1, 12) {real, imag} */,
  {32'h41974e47, 32'h42849da7} /* (28, 1, 11) {real, imag} */,
  {32'hc2b2b54e, 32'hc26197d0} /* (28, 1, 10) {real, imag} */,
  {32'h4223836c, 32'hc2669cff} /* (28, 1, 9) {real, imag} */,
  {32'h41f20306, 32'h429e6c5a} /* (28, 1, 8) {real, imag} */,
  {32'hc2676a1b, 32'h42b09d02} /* (28, 1, 7) {real, imag} */,
  {32'hc10ba4d6, 32'hc332fd9c} /* (28, 1, 6) {real, imag} */,
  {32'hc3539d83, 32'h42f76442} /* (28, 1, 5) {real, imag} */,
  {32'h41fcee46, 32'hc29caf3e} /* (28, 1, 4) {real, imag} */,
  {32'hc29ca86c, 32'hc1666372} /* (28, 1, 3) {real, imag} */,
  {32'h438e691d, 32'hc45a6975} /* (28, 1, 2) {real, imag} */,
  {32'h437c1e36, 32'h44a45798} /* (28, 1, 1) {real, imag} */,
  {32'h4357346e, 32'h00000000} /* (28, 1, 0) {real, imag} */,
  {32'h439e1560, 32'hc450d1c3} /* (28, 0, 31) {real, imag} */,
  {32'hc1a37d10, 32'h44287722} /* (28, 0, 30) {real, imag} */,
  {32'hc1f20efc, 32'hc29f58e8} /* (28, 0, 29) {real, imag} */,
  {32'h4249f8e6, 32'h4305261b} /* (28, 0, 28) {real, imag} */,
  {32'hc31fa41f, 32'hc11d6fb0} /* (28, 0, 27) {real, imag} */,
  {32'hc26d8f90, 32'hc246fe7e} /* (28, 0, 26) {real, imag} */,
  {32'h424d3fdb, 32'h41636396} /* (28, 0, 25) {real, imag} */,
  {32'h40413740, 32'h429ce1f0} /* (28, 0, 24) {real, imag} */,
  {32'hc0cb0448, 32'hc26eb256} /* (28, 0, 23) {real, imag} */,
  {32'h42077988, 32'h42328fa9} /* (28, 0, 22) {real, imag} */,
  {32'hc2aaecf2, 32'hc1cb98b8} /* (28, 0, 21) {real, imag} */,
  {32'h425dabb8, 32'h3fd1ee48} /* (28, 0, 20) {real, imag} */,
  {32'hc164ac54, 32'hc0659cd0} /* (28, 0, 19) {real, imag} */,
  {32'h41ca6c55, 32'h410bc596} /* (28, 0, 18) {real, imag} */,
  {32'h40ba24d0, 32'hc224ab08} /* (28, 0, 17) {real, imag} */,
  {32'h40b4754c, 32'h00000000} /* (28, 0, 16) {real, imag} */,
  {32'h40ba24d0, 32'h4224ab08} /* (28, 0, 15) {real, imag} */,
  {32'h41ca6c55, 32'hc10bc596} /* (28, 0, 14) {real, imag} */,
  {32'hc164ac54, 32'h40659cd0} /* (28, 0, 13) {real, imag} */,
  {32'h425dabb8, 32'hbfd1ee48} /* (28, 0, 12) {real, imag} */,
  {32'hc2aaecf2, 32'h41cb98b8} /* (28, 0, 11) {real, imag} */,
  {32'h42077988, 32'hc2328fa9} /* (28, 0, 10) {real, imag} */,
  {32'hc0cb0448, 32'h426eb256} /* (28, 0, 9) {real, imag} */,
  {32'h40413740, 32'hc29ce1f0} /* (28, 0, 8) {real, imag} */,
  {32'h424d3fdb, 32'hc1636396} /* (28, 0, 7) {real, imag} */,
  {32'hc26d8f90, 32'h4246fe7e} /* (28, 0, 6) {real, imag} */,
  {32'hc31fa41f, 32'h411d6fb0} /* (28, 0, 5) {real, imag} */,
  {32'h4249f8e6, 32'hc305261b} /* (28, 0, 4) {real, imag} */,
  {32'hc1f20efc, 32'h429f58e8} /* (28, 0, 3) {real, imag} */,
  {32'hc1a37d10, 32'hc4287722} /* (28, 0, 2) {real, imag} */,
  {32'h439e1560, 32'h4450d1c3} /* (28, 0, 1) {real, imag} */,
  {32'h41b11a40, 32'h00000000} /* (28, 0, 0) {real, imag} */,
  {32'h431b5c29, 32'hc2752780} /* (27, 31, 31) {real, imag} */,
  {32'hc390b6d6, 32'h43d6fd1b} /* (27, 31, 30) {real, imag} */,
  {32'hc3182dd0, 32'hc0847204} /* (27, 31, 29) {real, imag} */,
  {32'h430529ec, 32'h433cb236} /* (27, 31, 28) {real, imag} */,
  {32'hc2e7a235, 32'h4243f234} /* (27, 31, 27) {real, imag} */,
  {32'h42386360, 32'hc1da9e7d} /* (27, 31, 26) {real, imag} */,
  {32'h4090ea78, 32'h42825b28} /* (27, 31, 25) {real, imag} */,
  {32'h40615340, 32'h42579078} /* (27, 31, 24) {real, imag} */,
  {32'hc21ce11e, 32'h422e3d53} /* (27, 31, 23) {real, imag} */,
  {32'hc2a7cd1c, 32'hc28987e8} /* (27, 31, 22) {real, imag} */,
  {32'hc2439bb6, 32'hc1bf1dae} /* (27, 31, 21) {real, imag} */,
  {32'hc2a44412, 32'h414dbff0} /* (27, 31, 20) {real, imag} */,
  {32'h3de4ec00, 32'h3e856da0} /* (27, 31, 19) {real, imag} */,
  {32'h4146da00, 32'hc171012a} /* (27, 31, 18) {real, imag} */,
  {32'h41197e08, 32'hc2ad5b7b} /* (27, 31, 17) {real, imag} */,
  {32'h4253aaa8, 32'h00000000} /* (27, 31, 16) {real, imag} */,
  {32'h41197e08, 32'h42ad5b7b} /* (27, 31, 15) {real, imag} */,
  {32'h4146da00, 32'h4171012a} /* (27, 31, 14) {real, imag} */,
  {32'h3de4ec00, 32'hbe856da0} /* (27, 31, 13) {real, imag} */,
  {32'hc2a44412, 32'hc14dbff0} /* (27, 31, 12) {real, imag} */,
  {32'hc2439bb6, 32'h41bf1dae} /* (27, 31, 11) {real, imag} */,
  {32'hc2a7cd1c, 32'h428987e8} /* (27, 31, 10) {real, imag} */,
  {32'hc21ce11e, 32'hc22e3d53} /* (27, 31, 9) {real, imag} */,
  {32'h40615340, 32'hc2579078} /* (27, 31, 8) {real, imag} */,
  {32'h4090ea78, 32'hc2825b28} /* (27, 31, 7) {real, imag} */,
  {32'h42386360, 32'h41da9e7d} /* (27, 31, 6) {real, imag} */,
  {32'hc2e7a235, 32'hc243f234} /* (27, 31, 5) {real, imag} */,
  {32'h430529ec, 32'hc33cb236} /* (27, 31, 4) {real, imag} */,
  {32'hc3182dd0, 32'h40847204} /* (27, 31, 3) {real, imag} */,
  {32'hc390b6d6, 32'hc3d6fd1b} /* (27, 31, 2) {real, imag} */,
  {32'h431b5c29, 32'h42752780} /* (27, 31, 1) {real, imag} */,
  {32'hc42613e8, 32'h00000000} /* (27, 31, 0) {real, imag} */,
  {32'h44101014, 32'hc1b2d720} /* (27, 30, 31) {real, imag} */,
  {32'hc4266210, 32'h43c6820e} /* (27, 30, 30) {real, imag} */,
  {32'hc31dba3b, 32'hc1ab0602} /* (27, 30, 29) {real, imag} */,
  {32'h431e913f, 32'h433c6807} /* (27, 30, 28) {real, imag} */,
  {32'hc38bb51f, 32'h423e86b2} /* (27, 30, 27) {real, imag} */,
  {32'h4270c5e6, 32'h40b3e3c0} /* (27, 30, 26) {real, imag} */,
  {32'h429d7e38, 32'hc23f3094} /* (27, 30, 25) {real, imag} */,
  {32'hc16eff44, 32'h405e45f0} /* (27, 30, 24) {real, imag} */,
  {32'h41635950, 32'hc189f4cf} /* (27, 30, 23) {real, imag} */,
  {32'hc13dc20a, 32'hc2753e21} /* (27, 30, 22) {real, imag} */,
  {32'hc23fdecf, 32'hc24b4e86} /* (27, 30, 21) {real, imag} */,
  {32'hc3288604, 32'hc162992a} /* (27, 30, 20) {real, imag} */,
  {32'h4288b7d0, 32'h425f0373} /* (27, 30, 19) {real, imag} */,
  {32'h428ea969, 32'hc01d9680} /* (27, 30, 18) {real, imag} */,
  {32'h4200efa8, 32'hc19210d5} /* (27, 30, 17) {real, imag} */,
  {32'hc2c3eff6, 32'h00000000} /* (27, 30, 16) {real, imag} */,
  {32'h4200efa8, 32'h419210d5} /* (27, 30, 15) {real, imag} */,
  {32'h428ea969, 32'h401d9680} /* (27, 30, 14) {real, imag} */,
  {32'h4288b7d0, 32'hc25f0373} /* (27, 30, 13) {real, imag} */,
  {32'hc3288604, 32'h4162992a} /* (27, 30, 12) {real, imag} */,
  {32'hc23fdecf, 32'h424b4e86} /* (27, 30, 11) {real, imag} */,
  {32'hc13dc20a, 32'h42753e21} /* (27, 30, 10) {real, imag} */,
  {32'h41635950, 32'h4189f4cf} /* (27, 30, 9) {real, imag} */,
  {32'hc16eff44, 32'hc05e45f0} /* (27, 30, 8) {real, imag} */,
  {32'h429d7e38, 32'h423f3094} /* (27, 30, 7) {real, imag} */,
  {32'h4270c5e6, 32'hc0b3e3c0} /* (27, 30, 6) {real, imag} */,
  {32'hc38bb51f, 32'hc23e86b2} /* (27, 30, 5) {real, imag} */,
  {32'h431e913f, 32'hc33c6807} /* (27, 30, 4) {real, imag} */,
  {32'hc31dba3b, 32'h41ab0602} /* (27, 30, 3) {real, imag} */,
  {32'hc4266210, 32'hc3c6820e} /* (27, 30, 2) {real, imag} */,
  {32'h44101014, 32'h41b2d720} /* (27, 30, 1) {real, imag} */,
  {32'hc40a8758, 32'h00000000} /* (27, 30, 0) {real, imag} */,
  {32'h4438fca0, 32'h43374734} /* (27, 29, 31) {real, imag} */,
  {32'hc444bec0, 32'h43813b20} /* (27, 29, 30) {real, imag} */,
  {32'hc2cd4312, 32'h406f73b0} /* (27, 29, 29) {real, imag} */,
  {32'h41f52a9e, 32'hbf0a4a80} /* (27, 29, 28) {real, imag} */,
  {32'hc3933f55, 32'h426b2aaf} /* (27, 29, 27) {real, imag} */,
  {32'hc293d2be, 32'hc24338c2} /* (27, 29, 26) {real, imag} */,
  {32'h42114325, 32'hc2c61461} /* (27, 29, 25) {real, imag} */,
  {32'h42e00add, 32'h41d2c9de} /* (27, 29, 24) {real, imag} */,
  {32'h4206843a, 32'hc2b6f9e4} /* (27, 29, 23) {real, imag} */,
  {32'h4128aa08, 32'hc0d10a3c} /* (27, 29, 22) {real, imag} */,
  {32'hc200058f, 32'h4273f807} /* (27, 29, 21) {real, imag} */,
  {32'h413b67e4, 32'h424071f0} /* (27, 29, 20) {real, imag} */,
  {32'h4203e5b6, 32'h41fcf735} /* (27, 29, 19) {real, imag} */,
  {32'hc1cfd6f2, 32'hc0542ab0} /* (27, 29, 18) {real, imag} */,
  {32'h41d0d8f6, 32'hc20d5baf} /* (27, 29, 17) {real, imag} */,
  {32'hc2e16cc0, 32'h00000000} /* (27, 29, 16) {real, imag} */,
  {32'h41d0d8f6, 32'h420d5baf} /* (27, 29, 15) {real, imag} */,
  {32'hc1cfd6f2, 32'h40542ab0} /* (27, 29, 14) {real, imag} */,
  {32'h4203e5b6, 32'hc1fcf735} /* (27, 29, 13) {real, imag} */,
  {32'h413b67e4, 32'hc24071f0} /* (27, 29, 12) {real, imag} */,
  {32'hc200058f, 32'hc273f807} /* (27, 29, 11) {real, imag} */,
  {32'h4128aa08, 32'h40d10a3c} /* (27, 29, 10) {real, imag} */,
  {32'h4206843a, 32'h42b6f9e4} /* (27, 29, 9) {real, imag} */,
  {32'h42e00add, 32'hc1d2c9de} /* (27, 29, 8) {real, imag} */,
  {32'h42114325, 32'h42c61461} /* (27, 29, 7) {real, imag} */,
  {32'hc293d2be, 32'h424338c2} /* (27, 29, 6) {real, imag} */,
  {32'hc3933f55, 32'hc26b2aaf} /* (27, 29, 5) {real, imag} */,
  {32'h41f52a9e, 32'h3f0a4a80} /* (27, 29, 4) {real, imag} */,
  {32'hc2cd4312, 32'hc06f73b0} /* (27, 29, 3) {real, imag} */,
  {32'hc444bec0, 32'hc3813b20} /* (27, 29, 2) {real, imag} */,
  {32'h4438fca0, 32'hc3374734} /* (27, 29, 1) {real, imag} */,
  {32'hc3d96505, 32'h00000000} /* (27, 29, 0) {real, imag} */,
  {32'h44458346, 32'h43a2976d} /* (27, 28, 31) {real, imag} */,
  {32'hc44b13d2, 32'h4315d25c} /* (27, 28, 30) {real, imag} */,
  {32'hbef6c880, 32'hc26d230e} /* (27, 28, 29) {real, imag} */,
  {32'h43189c69, 32'hc1fb3ebf} /* (27, 28, 28) {real, imag} */,
  {32'hc36fb0c8, 32'h424531b5} /* (27, 28, 27) {real, imag} */,
  {32'h4253e553, 32'hc2a5085a} /* (27, 28, 26) {real, imag} */,
  {32'h42664564, 32'hc19a8608} /* (27, 28, 25) {real, imag} */,
  {32'hc2a38535, 32'h431bd6fc} /* (27, 28, 24) {real, imag} */,
  {32'hc30fa2a0, 32'hc24fee27} /* (27, 28, 23) {real, imag} */,
  {32'hc333f676, 32'hc107c9ca} /* (27, 28, 22) {real, imag} */,
  {32'h42d10b16, 32'h428a9822} /* (27, 28, 21) {real, imag} */,
  {32'h4283d59b, 32'hc2b8820d} /* (27, 28, 20) {real, imag} */,
  {32'h40982d60, 32'hc24f7bf2} /* (27, 28, 19) {real, imag} */,
  {32'h42a76e47, 32'h429378ae} /* (27, 28, 18) {real, imag} */,
  {32'h4240ecf4, 32'h41cf3d7a} /* (27, 28, 17) {real, imag} */,
  {32'hc1edd827, 32'h00000000} /* (27, 28, 16) {real, imag} */,
  {32'h4240ecf4, 32'hc1cf3d7a} /* (27, 28, 15) {real, imag} */,
  {32'h42a76e47, 32'hc29378ae} /* (27, 28, 14) {real, imag} */,
  {32'h40982d60, 32'h424f7bf2} /* (27, 28, 13) {real, imag} */,
  {32'h4283d59b, 32'h42b8820d} /* (27, 28, 12) {real, imag} */,
  {32'h42d10b16, 32'hc28a9822} /* (27, 28, 11) {real, imag} */,
  {32'hc333f676, 32'h4107c9ca} /* (27, 28, 10) {real, imag} */,
  {32'hc30fa2a0, 32'h424fee27} /* (27, 28, 9) {real, imag} */,
  {32'hc2a38535, 32'hc31bd6fc} /* (27, 28, 8) {real, imag} */,
  {32'h42664564, 32'h419a8608} /* (27, 28, 7) {real, imag} */,
  {32'h4253e553, 32'h42a5085a} /* (27, 28, 6) {real, imag} */,
  {32'hc36fb0c8, 32'hc24531b5} /* (27, 28, 5) {real, imag} */,
  {32'h43189c69, 32'h41fb3ebf} /* (27, 28, 4) {real, imag} */,
  {32'hbef6c880, 32'h426d230e} /* (27, 28, 3) {real, imag} */,
  {32'hc44b13d2, 32'hc315d25c} /* (27, 28, 2) {real, imag} */,
  {32'h44458346, 32'hc3a2976d} /* (27, 28, 1) {real, imag} */,
  {32'hc3b696f0, 32'h00000000} /* (27, 28, 0) {real, imag} */,
  {32'h443ecbc7, 32'h436d7f8e} /* (27, 27, 31) {real, imag} */,
  {32'hc451bf72, 32'h431e9910} /* (27, 27, 30) {real, imag} */,
  {32'h40364000, 32'hc2624108} /* (27, 27, 29) {real, imag} */,
  {32'hc107c915, 32'hc2fbafde} /* (27, 27, 28) {real, imag} */,
  {32'hc307925c, 32'h4371054c} /* (27, 27, 27) {real, imag} */,
  {32'h41c56996, 32'hc282c06d} /* (27, 27, 26) {real, imag} */,
  {32'h42be360e, 32'hc20effe4} /* (27, 27, 25) {real, imag} */,
  {32'hc269a326, 32'h42ce4618} /* (27, 27, 24) {real, imag} */,
  {32'hc2129415, 32'hc207402c} /* (27, 27, 23) {real, imag} */,
  {32'h4128d8ac, 32'hc1224d8c} /* (27, 27, 22) {real, imag} */,
  {32'h40ed2160, 32'h424ab3b1} /* (27, 27, 21) {real, imag} */,
  {32'h41c5aeb9, 32'hc189b90c} /* (27, 27, 20) {real, imag} */,
  {32'hc1a99ec2, 32'h414d3620} /* (27, 27, 19) {real, imag} */,
  {32'h41ae3902, 32'h426f4c1c} /* (27, 27, 18) {real, imag} */,
  {32'h41c3e826, 32'hc045c5d0} /* (27, 27, 17) {real, imag} */,
  {32'hc12cc226, 32'h00000000} /* (27, 27, 16) {real, imag} */,
  {32'h41c3e826, 32'h4045c5d0} /* (27, 27, 15) {real, imag} */,
  {32'h41ae3902, 32'hc26f4c1c} /* (27, 27, 14) {real, imag} */,
  {32'hc1a99ec2, 32'hc14d3620} /* (27, 27, 13) {real, imag} */,
  {32'h41c5aeb9, 32'h4189b90c} /* (27, 27, 12) {real, imag} */,
  {32'h40ed2160, 32'hc24ab3b1} /* (27, 27, 11) {real, imag} */,
  {32'h4128d8ac, 32'h41224d8c} /* (27, 27, 10) {real, imag} */,
  {32'hc2129415, 32'h4207402c} /* (27, 27, 9) {real, imag} */,
  {32'hc269a326, 32'hc2ce4618} /* (27, 27, 8) {real, imag} */,
  {32'h42be360e, 32'h420effe4} /* (27, 27, 7) {real, imag} */,
  {32'h41c56996, 32'h4282c06d} /* (27, 27, 6) {real, imag} */,
  {32'hc307925c, 32'hc371054c} /* (27, 27, 5) {real, imag} */,
  {32'hc107c915, 32'h42fbafde} /* (27, 27, 4) {real, imag} */,
  {32'h40364000, 32'h42624108} /* (27, 27, 3) {real, imag} */,
  {32'hc451bf72, 32'hc31e9910} /* (27, 27, 2) {real, imag} */,
  {32'h443ecbc7, 32'hc36d7f8e} /* (27, 27, 1) {real, imag} */,
  {32'hc3b3e658, 32'h00000000} /* (27, 27, 0) {real, imag} */,
  {32'h443c202d, 32'h4302224c} /* (27, 26, 31) {real, imag} */,
  {32'hc4551e0a, 32'h43618e23} /* (27, 26, 30) {real, imag} */,
  {32'h42675408, 32'hc21df60d} /* (27, 26, 29) {real, imag} */,
  {32'h430e4b0e, 32'hc2a68b03} /* (27, 26, 28) {real, imag} */,
  {32'hc2a5f138, 32'h4325880e} /* (27, 26, 27) {real, imag} */,
  {32'hc19d0f9c, 32'hc24a083e} /* (27, 26, 26) {real, imag} */,
  {32'h41a63ea8, 32'hc262f67e} /* (27, 26, 25) {real, imag} */,
  {32'hc1fa0d2c, 32'h42bbff0c} /* (27, 26, 24) {real, imag} */,
  {32'hc29d20a8, 32'h41344078} /* (27, 26, 23) {real, imag} */,
  {32'h4233d6b1, 32'hc20a9f38} /* (27, 26, 22) {real, imag} */,
  {32'hc28c78b0, 32'hc1c1a44e} /* (27, 26, 21) {real, imag} */,
  {32'h421f4fbe, 32'h428ea5a2} /* (27, 26, 20) {real, imag} */,
  {32'hc29f9570, 32'hc2933e89} /* (27, 26, 19) {real, imag} */,
  {32'h41c4ffc6, 32'h4266efdc} /* (27, 26, 18) {real, imag} */,
  {32'hc26cff77, 32'hc14601a8} /* (27, 26, 17) {real, imag} */,
  {32'hc0a35520, 32'h00000000} /* (27, 26, 16) {real, imag} */,
  {32'hc26cff77, 32'h414601a8} /* (27, 26, 15) {real, imag} */,
  {32'h41c4ffc6, 32'hc266efdc} /* (27, 26, 14) {real, imag} */,
  {32'hc29f9570, 32'h42933e89} /* (27, 26, 13) {real, imag} */,
  {32'h421f4fbe, 32'hc28ea5a2} /* (27, 26, 12) {real, imag} */,
  {32'hc28c78b0, 32'h41c1a44e} /* (27, 26, 11) {real, imag} */,
  {32'h4233d6b1, 32'h420a9f38} /* (27, 26, 10) {real, imag} */,
  {32'hc29d20a8, 32'hc1344078} /* (27, 26, 9) {real, imag} */,
  {32'hc1fa0d2c, 32'hc2bbff0c} /* (27, 26, 8) {real, imag} */,
  {32'h41a63ea8, 32'h4262f67e} /* (27, 26, 7) {real, imag} */,
  {32'hc19d0f9c, 32'h424a083e} /* (27, 26, 6) {real, imag} */,
  {32'hc2a5f138, 32'hc325880e} /* (27, 26, 5) {real, imag} */,
  {32'h430e4b0e, 32'h42a68b03} /* (27, 26, 4) {real, imag} */,
  {32'h42675408, 32'h421df60d} /* (27, 26, 3) {real, imag} */,
  {32'hc4551e0a, 32'hc3618e23} /* (27, 26, 2) {real, imag} */,
  {32'h443c202d, 32'hc302224c} /* (27, 26, 1) {real, imag} */,
  {32'hc4020968, 32'h00000000} /* (27, 26, 0) {real, imag} */,
  {32'h440c8318, 32'h42e5e564} /* (27, 25, 31) {real, imag} */,
  {32'hc44bb554, 32'h43655dc7} /* (27, 25, 30) {real, imag} */,
  {32'hc24542ec, 32'hc309c92e} /* (27, 25, 29) {real, imag} */,
  {32'h436ccc7d, 32'hc2624630} /* (27, 25, 28) {real, imag} */,
  {32'hc2b11f5e, 32'h41b8bf1c} /* (27, 25, 27) {real, imag} */,
  {32'hc2e77cad, 32'h42418716} /* (27, 25, 26) {real, imag} */,
  {32'hc19fbc3e, 32'hc305ee10} /* (27, 25, 25) {real, imag} */,
  {32'h400a9438, 32'h3e832740} /* (27, 25, 24) {real, imag} */,
  {32'hc2ed6a85, 32'h41f10e38} /* (27, 25, 23) {real, imag} */,
  {32'hc1dff177, 32'h40525e40} /* (27, 25, 22) {real, imag} */,
  {32'hc2e4ed1f, 32'h41f851c6} /* (27, 25, 21) {real, imag} */,
  {32'h42ed8bc9, 32'hc2892a5e} /* (27, 25, 20) {real, imag} */,
  {32'hc1864149, 32'hc15a1cd5} /* (27, 25, 19) {real, imag} */,
  {32'hc24b87cc, 32'hc253b3a2} /* (27, 25, 18) {real, imag} */,
  {32'h421501ea, 32'h410c35b4} /* (27, 25, 17) {real, imag} */,
  {32'h41b45679, 32'h00000000} /* (27, 25, 16) {real, imag} */,
  {32'h421501ea, 32'hc10c35b4} /* (27, 25, 15) {real, imag} */,
  {32'hc24b87cc, 32'h4253b3a2} /* (27, 25, 14) {real, imag} */,
  {32'hc1864149, 32'h415a1cd5} /* (27, 25, 13) {real, imag} */,
  {32'h42ed8bc9, 32'h42892a5e} /* (27, 25, 12) {real, imag} */,
  {32'hc2e4ed1f, 32'hc1f851c6} /* (27, 25, 11) {real, imag} */,
  {32'hc1dff177, 32'hc0525e40} /* (27, 25, 10) {real, imag} */,
  {32'hc2ed6a85, 32'hc1f10e38} /* (27, 25, 9) {real, imag} */,
  {32'h400a9438, 32'hbe832740} /* (27, 25, 8) {real, imag} */,
  {32'hc19fbc3e, 32'h4305ee10} /* (27, 25, 7) {real, imag} */,
  {32'hc2e77cad, 32'hc2418716} /* (27, 25, 6) {real, imag} */,
  {32'hc2b11f5e, 32'hc1b8bf1c} /* (27, 25, 5) {real, imag} */,
  {32'h436ccc7d, 32'h42624630} /* (27, 25, 4) {real, imag} */,
  {32'hc24542ec, 32'h4309c92e} /* (27, 25, 3) {real, imag} */,
  {32'hc44bb554, 32'hc3655dc7} /* (27, 25, 2) {real, imag} */,
  {32'h440c8318, 32'hc2e5e564} /* (27, 25, 1) {real, imag} */,
  {32'hc3b2d5ac, 32'h00000000} /* (27, 25, 0) {real, imag} */,
  {32'h44115f2b, 32'hc1041b34} /* (27, 24, 31) {real, imag} */,
  {32'hc450b2b9, 32'h4306328c} /* (27, 24, 30) {real, imag} */,
  {32'hc21cb9ab, 32'hc33b4fb5} /* (27, 24, 29) {real, imag} */,
  {32'h435732c0, 32'hc287aff0} /* (27, 24, 28) {real, imag} */,
  {32'hc2d8ccff, 32'h43398d5b} /* (27, 24, 27) {real, imag} */,
  {32'hc257f6c7, 32'h43055348} /* (27, 24, 26) {real, imag} */,
  {32'h42544be0, 32'hc33d54ba} /* (27, 24, 25) {real, imag} */,
  {32'hc1775a00, 32'h43243988} /* (27, 24, 24) {real, imag} */,
  {32'hc2de0592, 32'hc203cd77} /* (27, 24, 23) {real, imag} */,
  {32'h423c9ff9, 32'h42cde882} /* (27, 24, 22) {real, imag} */,
  {32'h426faec5, 32'h4212d88e} /* (27, 24, 21) {real, imag} */,
  {32'h42723ae8, 32'hbfef8140} /* (27, 24, 20) {real, imag} */,
  {32'hc29b0795, 32'h42a688c0} /* (27, 24, 19) {real, imag} */,
  {32'hc2552906, 32'h41683274} /* (27, 24, 18) {real, imag} */,
  {32'h42548ffe, 32'hc2aec486} /* (27, 24, 17) {real, imag} */,
  {32'hc1a4d401, 32'h00000000} /* (27, 24, 16) {real, imag} */,
  {32'h42548ffe, 32'h42aec486} /* (27, 24, 15) {real, imag} */,
  {32'hc2552906, 32'hc1683274} /* (27, 24, 14) {real, imag} */,
  {32'hc29b0795, 32'hc2a688c0} /* (27, 24, 13) {real, imag} */,
  {32'h42723ae8, 32'h3fef8140} /* (27, 24, 12) {real, imag} */,
  {32'h426faec5, 32'hc212d88e} /* (27, 24, 11) {real, imag} */,
  {32'h423c9ff9, 32'hc2cde882} /* (27, 24, 10) {real, imag} */,
  {32'hc2de0592, 32'h4203cd77} /* (27, 24, 9) {real, imag} */,
  {32'hc1775a00, 32'hc3243988} /* (27, 24, 8) {real, imag} */,
  {32'h42544be0, 32'h433d54ba} /* (27, 24, 7) {real, imag} */,
  {32'hc257f6c7, 32'hc3055348} /* (27, 24, 6) {real, imag} */,
  {32'hc2d8ccff, 32'hc3398d5b} /* (27, 24, 5) {real, imag} */,
  {32'h435732c0, 32'h4287aff0} /* (27, 24, 4) {real, imag} */,
  {32'hc21cb9ab, 32'h433b4fb5} /* (27, 24, 3) {real, imag} */,
  {32'hc450b2b9, 32'hc306328c} /* (27, 24, 2) {real, imag} */,
  {32'h44115f2b, 32'h41041b34} /* (27, 24, 1) {real, imag} */,
  {32'hc26dc6b2, 32'h00000000} /* (27, 24, 0) {real, imag} */,
  {32'h44033fd0, 32'hc1bbecfa} /* (27, 23, 31) {real, imag} */,
  {32'hc440b5d4, 32'h423d979e} /* (27, 23, 30) {real, imag} */,
  {32'h4220c324, 32'hc320fd98} /* (27, 23, 29) {real, imag} */,
  {32'h4320d34d, 32'hc27da526} /* (27, 23, 28) {real, imag} */,
  {32'hc34daaaf, 32'h432b9236} /* (27, 23, 27) {real, imag} */,
  {32'h415f057c, 32'h42d3ef1a} /* (27, 23, 26) {real, imag} */,
  {32'h425ffb8e, 32'hc2db164a} /* (27, 23, 25) {real, imag} */,
  {32'hc1c956f5, 32'hc12862d4} /* (27, 23, 24) {real, imag} */,
  {32'hc2e52675, 32'hc1f6536c} /* (27, 23, 23) {real, imag} */,
  {32'h423b855c, 32'h424e45fc} /* (27, 23, 22) {real, imag} */,
  {32'hc23a9ee4, 32'h42a79cda} /* (27, 23, 21) {real, imag} */,
  {32'h423c8156, 32'hc22baccc} /* (27, 23, 20) {real, imag} */,
  {32'h42a077f9, 32'h42129754} /* (27, 23, 19) {real, imag} */,
  {32'hc01bb740, 32'hc24948f0} /* (27, 23, 18) {real, imag} */,
  {32'h41e69cf6, 32'hc2976c14} /* (27, 23, 17) {real, imag} */,
  {32'h4247cde3, 32'h00000000} /* (27, 23, 16) {real, imag} */,
  {32'h41e69cf6, 32'h42976c14} /* (27, 23, 15) {real, imag} */,
  {32'hc01bb740, 32'h424948f0} /* (27, 23, 14) {real, imag} */,
  {32'h42a077f9, 32'hc2129754} /* (27, 23, 13) {real, imag} */,
  {32'h423c8156, 32'h422baccc} /* (27, 23, 12) {real, imag} */,
  {32'hc23a9ee4, 32'hc2a79cda} /* (27, 23, 11) {real, imag} */,
  {32'h423b855c, 32'hc24e45fc} /* (27, 23, 10) {real, imag} */,
  {32'hc2e52675, 32'h41f6536c} /* (27, 23, 9) {real, imag} */,
  {32'hc1c956f5, 32'h412862d4} /* (27, 23, 8) {real, imag} */,
  {32'h425ffb8e, 32'h42db164a} /* (27, 23, 7) {real, imag} */,
  {32'h415f057c, 32'hc2d3ef1a} /* (27, 23, 6) {real, imag} */,
  {32'hc34daaaf, 32'hc32b9236} /* (27, 23, 5) {real, imag} */,
  {32'h4320d34d, 32'h427da526} /* (27, 23, 4) {real, imag} */,
  {32'h4220c324, 32'h4320fd98} /* (27, 23, 3) {real, imag} */,
  {32'hc440b5d4, 32'hc23d979e} /* (27, 23, 2) {real, imag} */,
  {32'h44033fd0, 32'h41bbecfa} /* (27, 23, 1) {real, imag} */,
  {32'h4367073b, 32'h00000000} /* (27, 23, 0) {real, imag} */,
  {32'h43c97523, 32'h430f1908} /* (27, 22, 31) {real, imag} */,
  {32'hc3a9a31c, 32'hc0040440} /* (27, 22, 30) {real, imag} */,
  {32'h3f966740, 32'hc2481836} /* (27, 22, 29) {real, imag} */,
  {32'h4290917c, 32'hc2074fe4} /* (27, 22, 28) {real, imag} */,
  {32'hc2ea90d2, 32'h42b7692a} /* (27, 22, 27) {real, imag} */,
  {32'h42333042, 32'h42097f44} /* (27, 22, 26) {real, imag} */,
  {32'hc19fffec, 32'h418ad7ad} /* (27, 22, 25) {real, imag} */,
  {32'hc293aff5, 32'hc26ad622} /* (27, 22, 24) {real, imag} */,
  {32'h42931156, 32'h4250f48c} /* (27, 22, 23) {real, imag} */,
  {32'h424f8a02, 32'h4049428c} /* (27, 22, 22) {real, imag} */,
  {32'h412863ae, 32'h41f24cc3} /* (27, 22, 21) {real, imag} */,
  {32'h4207138c, 32'h412f8db7} /* (27, 22, 20) {real, imag} */,
  {32'h42126848, 32'hc209dec1} /* (27, 22, 19) {real, imag} */,
  {32'h41bd2696, 32'h42ccafa8} /* (27, 22, 18) {real, imag} */,
  {32'h3db3f7c0, 32'h41e57986} /* (27, 22, 17) {real, imag} */,
  {32'h4207f09f, 32'h00000000} /* (27, 22, 16) {real, imag} */,
  {32'h3db3f7c0, 32'hc1e57986} /* (27, 22, 15) {real, imag} */,
  {32'h41bd2696, 32'hc2ccafa8} /* (27, 22, 14) {real, imag} */,
  {32'h42126848, 32'h4209dec1} /* (27, 22, 13) {real, imag} */,
  {32'h4207138c, 32'hc12f8db7} /* (27, 22, 12) {real, imag} */,
  {32'h412863ae, 32'hc1f24cc3} /* (27, 22, 11) {real, imag} */,
  {32'h424f8a02, 32'hc049428c} /* (27, 22, 10) {real, imag} */,
  {32'h42931156, 32'hc250f48c} /* (27, 22, 9) {real, imag} */,
  {32'hc293aff5, 32'h426ad622} /* (27, 22, 8) {real, imag} */,
  {32'hc19fffec, 32'hc18ad7ad} /* (27, 22, 7) {real, imag} */,
  {32'h42333042, 32'hc2097f44} /* (27, 22, 6) {real, imag} */,
  {32'hc2ea90d2, 32'hc2b7692a} /* (27, 22, 5) {real, imag} */,
  {32'h4290917c, 32'h42074fe4} /* (27, 22, 4) {real, imag} */,
  {32'h3f966740, 32'h42481836} /* (27, 22, 3) {real, imag} */,
  {32'hc3a9a31c, 32'h40040440} /* (27, 22, 2) {real, imag} */,
  {32'h43c97523, 32'hc30f1908} /* (27, 22, 1) {real, imag} */,
  {32'h4330c978, 32'h00000000} /* (27, 22, 0) {real, imag} */,
  {32'hc32b0b03, 32'h435e448b} /* (27, 21, 31) {real, imag} */,
  {32'hc021eb80, 32'h40804a00} /* (27, 21, 30) {real, imag} */,
  {32'h41c1206c, 32'hc303d703} /* (27, 21, 29) {real, imag} */,
  {32'hc1f528e8, 32'h42eeaa96} /* (27, 21, 28) {real, imag} */,
  {32'hc16c418c, 32'h42a71cdb} /* (27, 21, 27) {real, imag} */,
  {32'hc1b1cc8a, 32'hc2001030} /* (27, 21, 26) {real, imag} */,
  {32'h42cdd7d2, 32'hc268c4e1} /* (27, 21, 25) {real, imag} */,
  {32'hc31c95c6, 32'h4188d5ca} /* (27, 21, 24) {real, imag} */,
  {32'hc1c3c797, 32'hc2f10f8a} /* (27, 21, 23) {real, imag} */,
  {32'h41fd20b4, 32'hc1c6cf20} /* (27, 21, 22) {real, imag} */,
  {32'h42df1ed0, 32'h40eb2aae} /* (27, 21, 21) {real, imag} */,
  {32'h41c6d03e, 32'h428aab0f} /* (27, 21, 20) {real, imag} */,
  {32'hc15d5f46, 32'hc10b3bc2} /* (27, 21, 19) {real, imag} */,
  {32'hc1ec2b30, 32'h419d20fd} /* (27, 21, 18) {real, imag} */,
  {32'h41c7ccbc, 32'h421b7f25} /* (27, 21, 17) {real, imag} */,
  {32'hc2bbcec9, 32'h00000000} /* (27, 21, 16) {real, imag} */,
  {32'h41c7ccbc, 32'hc21b7f25} /* (27, 21, 15) {real, imag} */,
  {32'hc1ec2b30, 32'hc19d20fd} /* (27, 21, 14) {real, imag} */,
  {32'hc15d5f46, 32'h410b3bc2} /* (27, 21, 13) {real, imag} */,
  {32'h41c6d03e, 32'hc28aab0f} /* (27, 21, 12) {real, imag} */,
  {32'h42df1ed0, 32'hc0eb2aae} /* (27, 21, 11) {real, imag} */,
  {32'h41fd20b4, 32'h41c6cf20} /* (27, 21, 10) {real, imag} */,
  {32'hc1c3c797, 32'h42f10f8a} /* (27, 21, 9) {real, imag} */,
  {32'hc31c95c6, 32'hc188d5ca} /* (27, 21, 8) {real, imag} */,
  {32'h42cdd7d2, 32'h4268c4e1} /* (27, 21, 7) {real, imag} */,
  {32'hc1b1cc8a, 32'h42001030} /* (27, 21, 6) {real, imag} */,
  {32'hc16c418c, 32'hc2a71cdb} /* (27, 21, 5) {real, imag} */,
  {32'hc1f528e8, 32'hc2eeaa96} /* (27, 21, 4) {real, imag} */,
  {32'h41c1206c, 32'h4303d703} /* (27, 21, 3) {real, imag} */,
  {32'hc021eb80, 32'hc0804a00} /* (27, 21, 2) {real, imag} */,
  {32'hc32b0b03, 32'hc35e448b} /* (27, 21, 1) {real, imag} */,
  {32'hc0dbbb00, 32'h00000000} /* (27, 21, 0) {real, imag} */,
  {32'hc4720e8f, 32'h4332cfc3} /* (27, 20, 31) {real, imag} */,
  {32'h43f65f8e, 32'hc2b5937c} /* (27, 20, 30) {real, imag} */,
  {32'hc1bc8ec7, 32'hc30390ce} /* (27, 20, 29) {real, imag} */,
  {32'h41c652e8, 32'h42109720} /* (27, 20, 28) {real, imag} */,
  {32'h428744c4, 32'hc29786cc} /* (27, 20, 27) {real, imag} */,
  {32'h419c2f36, 32'h407602e8} /* (27, 20, 26) {real, imag} */,
  {32'h42760385, 32'hc2e75346} /* (27, 20, 25) {real, imag} */,
  {32'hc26f2113, 32'hc1d79b8c} /* (27, 20, 24) {real, imag} */,
  {32'hc2ba39c2, 32'h41e4e314} /* (27, 20, 23) {real, imag} */,
  {32'hc22ab6cc, 32'h42ac13de} /* (27, 20, 22) {real, imag} */,
  {32'h42ab5ea1, 32'h4254057d} /* (27, 20, 21) {real, imag} */,
  {32'h423a0da4, 32'hc28d2d9c} /* (27, 20, 20) {real, imag} */,
  {32'hc23f47b6, 32'hc1440bb4} /* (27, 20, 19) {real, imag} */,
  {32'h422dfec4, 32'hc2339d65} /* (27, 20, 18) {real, imag} */,
  {32'hc247b529, 32'hc164e1e0} /* (27, 20, 17) {real, imag} */,
  {32'h4212f652, 32'h00000000} /* (27, 20, 16) {real, imag} */,
  {32'hc247b529, 32'h4164e1e0} /* (27, 20, 15) {real, imag} */,
  {32'h422dfec4, 32'h42339d65} /* (27, 20, 14) {real, imag} */,
  {32'hc23f47b6, 32'h41440bb4} /* (27, 20, 13) {real, imag} */,
  {32'h423a0da4, 32'h428d2d9c} /* (27, 20, 12) {real, imag} */,
  {32'h42ab5ea1, 32'hc254057d} /* (27, 20, 11) {real, imag} */,
  {32'hc22ab6cc, 32'hc2ac13de} /* (27, 20, 10) {real, imag} */,
  {32'hc2ba39c2, 32'hc1e4e314} /* (27, 20, 9) {real, imag} */,
  {32'hc26f2113, 32'h41d79b8c} /* (27, 20, 8) {real, imag} */,
  {32'h42760385, 32'h42e75346} /* (27, 20, 7) {real, imag} */,
  {32'h419c2f36, 32'hc07602e8} /* (27, 20, 6) {real, imag} */,
  {32'h428744c4, 32'h429786cc} /* (27, 20, 5) {real, imag} */,
  {32'h41c652e8, 32'hc2109720} /* (27, 20, 4) {real, imag} */,
  {32'hc1bc8ec7, 32'h430390ce} /* (27, 20, 3) {real, imag} */,
  {32'h43f65f8e, 32'h42b5937c} /* (27, 20, 2) {real, imag} */,
  {32'hc4720e8f, 32'hc332cfc3} /* (27, 20, 1) {real, imag} */,
  {32'hc40bb049, 32'h00000000} /* (27, 20, 0) {real, imag} */,
  {32'hc495f8ca, 32'h4373b1bd} /* (27, 19, 31) {real, imag} */,
  {32'h4418a2dc, 32'hc37631d0} /* (27, 19, 30) {real, imag} */,
  {32'h40bb89c0, 32'hc3002b68} /* (27, 19, 29) {real, imag} */,
  {32'hc1734244, 32'hc2116ff8} /* (27, 19, 28) {real, imag} */,
  {32'h43097302, 32'h4138134c} /* (27, 19, 27) {real, imag} */,
  {32'h42866972, 32'hc2877b67} /* (27, 19, 26) {real, imag} */,
  {32'hc19be5c6, 32'h4289df8e} /* (27, 19, 25) {real, imag} */,
  {32'h41fd1f0a, 32'h42075912} /* (27, 19, 24) {real, imag} */,
  {32'h42c3cf6d, 32'h4199d49e} /* (27, 19, 23) {real, imag} */,
  {32'h42b78f98, 32'h4208db76} /* (27, 19, 22) {real, imag} */,
  {32'h428845fc, 32'h4274772d} /* (27, 19, 21) {real, imag} */,
  {32'hc2aa9182, 32'h42b60b03} /* (27, 19, 20) {real, imag} */,
  {32'h40e69864, 32'h42bf7a63} /* (27, 19, 19) {real, imag} */,
  {32'hc262fe99, 32'hc1cc083d} /* (27, 19, 18) {real, imag} */,
  {32'h411ae7bb, 32'h41ae7dda} /* (27, 19, 17) {real, imag} */,
  {32'hc11c7744, 32'h00000000} /* (27, 19, 16) {real, imag} */,
  {32'h411ae7bb, 32'hc1ae7dda} /* (27, 19, 15) {real, imag} */,
  {32'hc262fe99, 32'h41cc083d} /* (27, 19, 14) {real, imag} */,
  {32'h40e69864, 32'hc2bf7a63} /* (27, 19, 13) {real, imag} */,
  {32'hc2aa9182, 32'hc2b60b03} /* (27, 19, 12) {real, imag} */,
  {32'h428845fc, 32'hc274772d} /* (27, 19, 11) {real, imag} */,
  {32'h42b78f98, 32'hc208db76} /* (27, 19, 10) {real, imag} */,
  {32'h42c3cf6d, 32'hc199d49e} /* (27, 19, 9) {real, imag} */,
  {32'h41fd1f0a, 32'hc2075912} /* (27, 19, 8) {real, imag} */,
  {32'hc19be5c6, 32'hc289df8e} /* (27, 19, 7) {real, imag} */,
  {32'h42866972, 32'h42877b67} /* (27, 19, 6) {real, imag} */,
  {32'h43097302, 32'hc138134c} /* (27, 19, 5) {real, imag} */,
  {32'hc1734244, 32'h42116ff8} /* (27, 19, 4) {real, imag} */,
  {32'h40bb89c0, 32'h43002b68} /* (27, 19, 3) {real, imag} */,
  {32'h4418a2dc, 32'h437631d0} /* (27, 19, 2) {real, imag} */,
  {32'hc495f8ca, 32'hc373b1bd} /* (27, 19, 1) {real, imag} */,
  {32'hc4267762, 32'h00000000} /* (27, 19, 0) {real, imag} */,
  {32'hc49dd857, 32'h43af8800} /* (27, 18, 31) {real, imag} */,
  {32'h443ee154, 32'hc3a1ab68} /* (27, 18, 30) {real, imag} */,
  {32'h42e20868, 32'hc1875a72} /* (27, 18, 29) {real, imag} */,
  {32'hc1a74160, 32'h431493d7} /* (27, 18, 28) {real, imag} */,
  {32'h4294f67b, 32'h42b451dc} /* (27, 18, 27) {real, imag} */,
  {32'hc0a747d8, 32'h420979e2} /* (27, 18, 26) {real, imag} */,
  {32'hc183f23d, 32'hc293833c} /* (27, 18, 25) {real, imag} */,
  {32'h4251680c, 32'h41cd9968} /* (27, 18, 24) {real, imag} */,
  {32'h421f9b96, 32'h40a44eaa} /* (27, 18, 23) {real, imag} */,
  {32'hc1b7f09d, 32'h3fea0680} /* (27, 18, 22) {real, imag} */,
  {32'hc263ef74, 32'h41962853} /* (27, 18, 21) {real, imag} */,
  {32'hc145455c, 32'hc2bc932f} /* (27, 18, 20) {real, imag} */,
  {32'hc214483e, 32'h41aa84f2} /* (27, 18, 19) {real, imag} */,
  {32'h42d6fa0e, 32'hc2731224} /* (27, 18, 18) {real, imag} */,
  {32'h42a84736, 32'hc10e85e2} /* (27, 18, 17) {real, imag} */,
  {32'hc21304dc, 32'h00000000} /* (27, 18, 16) {real, imag} */,
  {32'h42a84736, 32'h410e85e2} /* (27, 18, 15) {real, imag} */,
  {32'h42d6fa0e, 32'h42731224} /* (27, 18, 14) {real, imag} */,
  {32'hc214483e, 32'hc1aa84f2} /* (27, 18, 13) {real, imag} */,
  {32'hc145455c, 32'h42bc932f} /* (27, 18, 12) {real, imag} */,
  {32'hc263ef74, 32'hc1962853} /* (27, 18, 11) {real, imag} */,
  {32'hc1b7f09d, 32'hbfea0680} /* (27, 18, 10) {real, imag} */,
  {32'h421f9b96, 32'hc0a44eaa} /* (27, 18, 9) {real, imag} */,
  {32'h4251680c, 32'hc1cd9968} /* (27, 18, 8) {real, imag} */,
  {32'hc183f23d, 32'h4293833c} /* (27, 18, 7) {real, imag} */,
  {32'hc0a747d8, 32'hc20979e2} /* (27, 18, 6) {real, imag} */,
  {32'h4294f67b, 32'hc2b451dc} /* (27, 18, 5) {real, imag} */,
  {32'hc1a74160, 32'hc31493d7} /* (27, 18, 4) {real, imag} */,
  {32'h42e20868, 32'h41875a72} /* (27, 18, 3) {real, imag} */,
  {32'h443ee154, 32'h43a1ab68} /* (27, 18, 2) {real, imag} */,
  {32'hc49dd857, 32'hc3af8800} /* (27, 18, 1) {real, imag} */,
  {32'hc459088e, 32'h00000000} /* (27, 18, 0) {real, imag} */,
  {32'hc49fade5, 32'h43a721e4} /* (27, 17, 31) {real, imag} */,
  {32'h4440c880, 32'hc359a3e8} /* (27, 17, 30) {real, imag} */,
  {32'hbf997050, 32'hc2b2c3b2} /* (27, 17, 29) {real, imag} */,
  {32'h422e3055, 32'h436074bb} /* (27, 17, 28) {real, imag} */,
  {32'h433a738e, 32'hc28a56db} /* (27, 17, 27) {real, imag} */,
  {32'h42eea554, 32'h414a4812} /* (27, 17, 26) {real, imag} */,
  {32'h429052d7, 32'hc2ec9c77} /* (27, 17, 25) {real, imag} */,
  {32'h41c9e6b1, 32'hc113f388} /* (27, 17, 24) {real, imag} */,
  {32'h429d21d1, 32'h4210d7f5} /* (27, 17, 23) {real, imag} */,
  {32'h42411766, 32'h42f542d9} /* (27, 17, 22) {real, imag} */,
  {32'hc127d564, 32'hc2d1f185} /* (27, 17, 21) {real, imag} */,
  {32'h407f9190, 32'h42654b49} /* (27, 17, 20) {real, imag} */,
  {32'h41551f98, 32'h411a503c} /* (27, 17, 19) {real, imag} */,
  {32'hc21e9dee, 32'h424cfd74} /* (27, 17, 18) {real, imag} */,
  {32'hc0549ee0, 32'h42bb9f5a} /* (27, 17, 17) {real, imag} */,
  {32'hc21f134c, 32'h00000000} /* (27, 17, 16) {real, imag} */,
  {32'hc0549ee0, 32'hc2bb9f5a} /* (27, 17, 15) {real, imag} */,
  {32'hc21e9dee, 32'hc24cfd74} /* (27, 17, 14) {real, imag} */,
  {32'h41551f98, 32'hc11a503c} /* (27, 17, 13) {real, imag} */,
  {32'h407f9190, 32'hc2654b49} /* (27, 17, 12) {real, imag} */,
  {32'hc127d564, 32'h42d1f185} /* (27, 17, 11) {real, imag} */,
  {32'h42411766, 32'hc2f542d9} /* (27, 17, 10) {real, imag} */,
  {32'h429d21d1, 32'hc210d7f5} /* (27, 17, 9) {real, imag} */,
  {32'h41c9e6b1, 32'h4113f388} /* (27, 17, 8) {real, imag} */,
  {32'h429052d7, 32'h42ec9c77} /* (27, 17, 7) {real, imag} */,
  {32'h42eea554, 32'hc14a4812} /* (27, 17, 6) {real, imag} */,
  {32'h433a738e, 32'h428a56db} /* (27, 17, 5) {real, imag} */,
  {32'h422e3055, 32'hc36074bb} /* (27, 17, 4) {real, imag} */,
  {32'hbf997050, 32'h42b2c3b2} /* (27, 17, 3) {real, imag} */,
  {32'h4440c880, 32'h4359a3e8} /* (27, 17, 2) {real, imag} */,
  {32'hc49fade5, 32'hc3a721e4} /* (27, 17, 1) {real, imag} */,
  {32'hc476fe8e, 32'h00000000} /* (27, 17, 0) {real, imag} */,
  {32'hc49ebafa, 32'h438d8580} /* (27, 16, 31) {real, imag} */,
  {32'h442c113c, 32'hc2eefd58} /* (27, 16, 30) {real, imag} */,
  {32'h4290fa18, 32'hc2b64edd} /* (27, 16, 29) {real, imag} */,
  {32'hc2ec243f, 32'h42c55686} /* (27, 16, 28) {real, imag} */,
  {32'h432ef188, 32'h41495b8c} /* (27, 16, 27) {real, imag} */,
  {32'h4267cd92, 32'h3f1ce550} /* (27, 16, 26) {real, imag} */,
  {32'h40219370, 32'hc236f3c3} /* (27, 16, 25) {real, imag} */,
  {32'h4283ea7f, 32'hc2635194} /* (27, 16, 24) {real, imag} */,
  {32'hc243c8dd, 32'hc113c867} /* (27, 16, 23) {real, imag} */,
  {32'hc2bc56fc, 32'hc280b1fa} /* (27, 16, 22) {real, imag} */,
  {32'h410db3aa, 32'hc2750cc8} /* (27, 16, 21) {real, imag} */,
  {32'h40c1868c, 32'hc1eeae29} /* (27, 16, 20) {real, imag} */,
  {32'hc175ec42, 32'hc1e47e2a} /* (27, 16, 19) {real, imag} */,
  {32'hc27b0712, 32'h40a4bb90} /* (27, 16, 18) {real, imag} */,
  {32'h420fd2be, 32'h42a8b736} /* (27, 16, 17) {real, imag} */,
  {32'hc1aba374, 32'h00000000} /* (27, 16, 16) {real, imag} */,
  {32'h420fd2be, 32'hc2a8b736} /* (27, 16, 15) {real, imag} */,
  {32'hc27b0712, 32'hc0a4bb90} /* (27, 16, 14) {real, imag} */,
  {32'hc175ec42, 32'h41e47e2a} /* (27, 16, 13) {real, imag} */,
  {32'h40c1868c, 32'h41eeae29} /* (27, 16, 12) {real, imag} */,
  {32'h410db3aa, 32'h42750cc8} /* (27, 16, 11) {real, imag} */,
  {32'hc2bc56fc, 32'h4280b1fa} /* (27, 16, 10) {real, imag} */,
  {32'hc243c8dd, 32'h4113c867} /* (27, 16, 9) {real, imag} */,
  {32'h4283ea7f, 32'h42635194} /* (27, 16, 8) {real, imag} */,
  {32'h40219370, 32'h4236f3c3} /* (27, 16, 7) {real, imag} */,
  {32'h4267cd92, 32'hbf1ce550} /* (27, 16, 6) {real, imag} */,
  {32'h432ef188, 32'hc1495b8c} /* (27, 16, 5) {real, imag} */,
  {32'hc2ec243f, 32'hc2c55686} /* (27, 16, 4) {real, imag} */,
  {32'h4290fa18, 32'h42b64edd} /* (27, 16, 3) {real, imag} */,
  {32'h442c113c, 32'h42eefd58} /* (27, 16, 2) {real, imag} */,
  {32'hc49ebafa, 32'hc38d8580} /* (27, 16, 1) {real, imag} */,
  {32'hc484ff20, 32'h00000000} /* (27, 16, 0) {real, imag} */,
  {32'hc48c422f, 32'h43923984} /* (27, 15, 31) {real, imag} */,
  {32'h4438228a, 32'hc2a87338} /* (27, 15, 30) {real, imag} */,
  {32'h4229f956, 32'hc24ed1dc} /* (27, 15, 29) {real, imag} */,
  {32'hc2c41b0c, 32'h42ec7ab2} /* (27, 15, 28) {real, imag} */,
  {32'h42a8ae8c, 32'hc2a9b10d} /* (27, 15, 27) {real, imag} */,
  {32'hc24c8681, 32'hc188a6a3} /* (27, 15, 26) {real, imag} */,
  {32'hc23c4f92, 32'h42b74e11} /* (27, 15, 25) {real, imag} */,
  {32'h42aa112a, 32'hc30adbf2} /* (27, 15, 24) {real, imag} */,
  {32'hc1ede169, 32'hc182cf66} /* (27, 15, 23) {real, imag} */,
  {32'hc27aa0da, 32'h42d8770b} /* (27, 15, 22) {real, imag} */,
  {32'h42185103, 32'hc21efd8e} /* (27, 15, 21) {real, imag} */,
  {32'h42271a25, 32'h3ec55d80} /* (27, 15, 20) {real, imag} */,
  {32'hbed17b40, 32'h4253f90f} /* (27, 15, 19) {real, imag} */,
  {32'h42692b96, 32'hc294b422} /* (27, 15, 18) {real, imag} */,
  {32'h42c3f64d, 32'hc210b9f1} /* (27, 15, 17) {real, imag} */,
  {32'hc2abfdd2, 32'h00000000} /* (27, 15, 16) {real, imag} */,
  {32'h42c3f64d, 32'h4210b9f1} /* (27, 15, 15) {real, imag} */,
  {32'h42692b96, 32'h4294b422} /* (27, 15, 14) {real, imag} */,
  {32'hbed17b40, 32'hc253f90f} /* (27, 15, 13) {real, imag} */,
  {32'h42271a25, 32'hbec55d80} /* (27, 15, 12) {real, imag} */,
  {32'h42185103, 32'h421efd8e} /* (27, 15, 11) {real, imag} */,
  {32'hc27aa0da, 32'hc2d8770b} /* (27, 15, 10) {real, imag} */,
  {32'hc1ede169, 32'h4182cf66} /* (27, 15, 9) {real, imag} */,
  {32'h42aa112a, 32'h430adbf2} /* (27, 15, 8) {real, imag} */,
  {32'hc23c4f92, 32'hc2b74e11} /* (27, 15, 7) {real, imag} */,
  {32'hc24c8681, 32'h4188a6a3} /* (27, 15, 6) {real, imag} */,
  {32'h42a8ae8c, 32'h42a9b10d} /* (27, 15, 5) {real, imag} */,
  {32'hc2c41b0c, 32'hc2ec7ab2} /* (27, 15, 4) {real, imag} */,
  {32'h4229f956, 32'h424ed1dc} /* (27, 15, 3) {real, imag} */,
  {32'h4438228a, 32'h42a87338} /* (27, 15, 2) {real, imag} */,
  {32'hc48c422f, 32'hc3923984} /* (27, 15, 1) {real, imag} */,
  {32'hc4988a5f, 32'h00000000} /* (27, 15, 0) {real, imag} */,
  {32'hc484f901, 32'h43a38156} /* (27, 14, 31) {real, imag} */,
  {32'h442d011c, 32'hc1ff6808} /* (27, 14, 30) {real, imag} */,
  {32'hc0c00c38, 32'h41245618} /* (27, 14, 29) {real, imag} */,
  {32'hc33457f8, 32'h42d626d3} /* (27, 14, 28) {real, imag} */,
  {32'h43359a28, 32'hc2e684a0} /* (27, 14, 27) {real, imag} */,
  {32'h429f129c, 32'hc1e19c3a} /* (27, 14, 26) {real, imag} */,
  {32'hc052f428, 32'h42779a88} /* (27, 14, 25) {real, imag} */,
  {32'h42613042, 32'hc1f41200} /* (27, 14, 24) {real, imag} */,
  {32'h42401c9c, 32'h418c32e0} /* (27, 14, 23) {real, imag} */,
  {32'h4198b283, 32'hc2a7b803} /* (27, 14, 22) {real, imag} */,
  {32'h43194f5d, 32'hc181d9cf} /* (27, 14, 21) {real, imag} */,
  {32'h429f620e, 32'hc2ae0141} /* (27, 14, 20) {real, imag} */,
  {32'hc0eccf74, 32'hc088c6a6} /* (27, 14, 19) {real, imag} */,
  {32'h4118c7b0, 32'hc1e936ef} /* (27, 14, 18) {real, imag} */,
  {32'hc0997220, 32'hc2242398} /* (27, 14, 17) {real, imag} */,
  {32'h41f944a0, 32'h00000000} /* (27, 14, 16) {real, imag} */,
  {32'hc0997220, 32'h42242398} /* (27, 14, 15) {real, imag} */,
  {32'h4118c7b0, 32'h41e936ef} /* (27, 14, 14) {real, imag} */,
  {32'hc0eccf74, 32'h4088c6a6} /* (27, 14, 13) {real, imag} */,
  {32'h429f620e, 32'h42ae0141} /* (27, 14, 12) {real, imag} */,
  {32'h43194f5d, 32'h4181d9cf} /* (27, 14, 11) {real, imag} */,
  {32'h4198b283, 32'h42a7b803} /* (27, 14, 10) {real, imag} */,
  {32'h42401c9c, 32'hc18c32e0} /* (27, 14, 9) {real, imag} */,
  {32'h42613042, 32'h41f41200} /* (27, 14, 8) {real, imag} */,
  {32'hc052f428, 32'hc2779a88} /* (27, 14, 7) {real, imag} */,
  {32'h429f129c, 32'h41e19c3a} /* (27, 14, 6) {real, imag} */,
  {32'h43359a28, 32'h42e684a0} /* (27, 14, 5) {real, imag} */,
  {32'hc33457f8, 32'hc2d626d3} /* (27, 14, 4) {real, imag} */,
  {32'hc0c00c38, 32'hc1245618} /* (27, 14, 3) {real, imag} */,
  {32'h442d011c, 32'h41ff6808} /* (27, 14, 2) {real, imag} */,
  {32'hc484f901, 32'hc3a38156} /* (27, 14, 1) {real, imag} */,
  {32'hc48f5b72, 32'h00000000} /* (27, 14, 0) {real, imag} */,
  {32'hc46b0098, 32'h43520d57} /* (27, 13, 31) {real, imag} */,
  {32'h440bd284, 32'hc2683660} /* (27, 13, 30) {real, imag} */,
  {32'hc26407dc, 32'h428a91c4} /* (27, 13, 29) {real, imag} */,
  {32'hc30258f6, 32'h42df06b6} /* (27, 13, 28) {real, imag} */,
  {32'h42faced8, 32'hc30b201c} /* (27, 13, 27) {real, imag} */,
  {32'h431adc25, 32'h4296c665} /* (27, 13, 26) {real, imag} */,
  {32'h426e4705, 32'hc0f2ab6c} /* (27, 13, 25) {real, imag} */,
  {32'h41f290c0, 32'h425447ac} /* (27, 13, 24) {real, imag} */,
  {32'h3eee2d00, 32'h42abc372} /* (27, 13, 23) {real, imag} */,
  {32'hc1dd1758, 32'hc02bbe08} /* (27, 13, 22) {real, imag} */,
  {32'h413b2848, 32'hc2d96eb6} /* (27, 13, 21) {real, imag} */,
  {32'h424a55cc, 32'h4183dfb0} /* (27, 13, 20) {real, imag} */,
  {32'hc1a1ddd3, 32'h4188027c} /* (27, 13, 19) {real, imag} */,
  {32'hc2317585, 32'hc199e16b} /* (27, 13, 18) {real, imag} */,
  {32'hc0fa7a56, 32'h4145fba3} /* (27, 13, 17) {real, imag} */,
  {32'h42f1454c, 32'h00000000} /* (27, 13, 16) {real, imag} */,
  {32'hc0fa7a56, 32'hc145fba3} /* (27, 13, 15) {real, imag} */,
  {32'hc2317585, 32'h4199e16b} /* (27, 13, 14) {real, imag} */,
  {32'hc1a1ddd3, 32'hc188027c} /* (27, 13, 13) {real, imag} */,
  {32'h424a55cc, 32'hc183dfb0} /* (27, 13, 12) {real, imag} */,
  {32'h413b2848, 32'h42d96eb6} /* (27, 13, 11) {real, imag} */,
  {32'hc1dd1758, 32'h402bbe08} /* (27, 13, 10) {real, imag} */,
  {32'h3eee2d00, 32'hc2abc372} /* (27, 13, 9) {real, imag} */,
  {32'h41f290c0, 32'hc25447ac} /* (27, 13, 8) {real, imag} */,
  {32'h426e4705, 32'h40f2ab6c} /* (27, 13, 7) {real, imag} */,
  {32'h431adc25, 32'hc296c665} /* (27, 13, 6) {real, imag} */,
  {32'h42faced8, 32'h430b201c} /* (27, 13, 5) {real, imag} */,
  {32'hc30258f6, 32'hc2df06b6} /* (27, 13, 4) {real, imag} */,
  {32'hc26407dc, 32'hc28a91c4} /* (27, 13, 3) {real, imag} */,
  {32'h440bd284, 32'h42683660} /* (27, 13, 2) {real, imag} */,
  {32'hc46b0098, 32'hc3520d57} /* (27, 13, 1) {real, imag} */,
  {32'hc4845779, 32'h00000000} /* (27, 13, 0) {real, imag} */,
  {32'hc44267a1, 32'h4371be91} /* (27, 12, 31) {real, imag} */,
  {32'h43d72910, 32'hc20b3ff0} /* (27, 12, 30) {real, imag} */,
  {32'hc04c9f28, 32'hc13fd0e8} /* (27, 12, 29) {real, imag} */,
  {32'hc20bca42, 32'h423d6d88} /* (27, 12, 28) {real, imag} */,
  {32'h41a832d7, 32'hc29f0b4c} /* (27, 12, 27) {real, imag} */,
  {32'hc1d7f8ca, 32'h42032e48} /* (27, 12, 26) {real, imag} */,
  {32'h422a1e8b, 32'hc1d2b916} /* (27, 12, 25) {real, imag} */,
  {32'h424a6759, 32'h41921604} /* (27, 12, 24) {real, imag} */,
  {32'h42ae0ffe, 32'hc1caed28} /* (27, 12, 23) {real, imag} */,
  {32'hc2c6f642, 32'h4327c0ac} /* (27, 12, 22) {real, imag} */,
  {32'h4232d6b2, 32'hc2078dbd} /* (27, 12, 21) {real, imag} */,
  {32'h42da0344, 32'hc26ce595} /* (27, 12, 20) {real, imag} */,
  {32'hc2890c85, 32'h41622a66} /* (27, 12, 19) {real, imag} */,
  {32'hc116692e, 32'hbd7e3800} /* (27, 12, 18) {real, imag} */,
  {32'h41d119f2, 32'hc1a249d8} /* (27, 12, 17) {real, imag} */,
  {32'hc2a7810b, 32'h00000000} /* (27, 12, 16) {real, imag} */,
  {32'h41d119f2, 32'h41a249d8} /* (27, 12, 15) {real, imag} */,
  {32'hc116692e, 32'h3d7e3800} /* (27, 12, 14) {real, imag} */,
  {32'hc2890c85, 32'hc1622a66} /* (27, 12, 13) {real, imag} */,
  {32'h42da0344, 32'h426ce595} /* (27, 12, 12) {real, imag} */,
  {32'h4232d6b2, 32'h42078dbd} /* (27, 12, 11) {real, imag} */,
  {32'hc2c6f642, 32'hc327c0ac} /* (27, 12, 10) {real, imag} */,
  {32'h42ae0ffe, 32'h41caed28} /* (27, 12, 9) {real, imag} */,
  {32'h424a6759, 32'hc1921604} /* (27, 12, 8) {real, imag} */,
  {32'h422a1e8b, 32'h41d2b916} /* (27, 12, 7) {real, imag} */,
  {32'hc1d7f8ca, 32'hc2032e48} /* (27, 12, 6) {real, imag} */,
  {32'h41a832d7, 32'h429f0b4c} /* (27, 12, 5) {real, imag} */,
  {32'hc20bca42, 32'hc23d6d88} /* (27, 12, 4) {real, imag} */,
  {32'hc04c9f28, 32'h413fd0e8} /* (27, 12, 3) {real, imag} */,
  {32'h43d72910, 32'h420b3ff0} /* (27, 12, 2) {real, imag} */,
  {32'hc44267a1, 32'hc371be91} /* (27, 12, 1) {real, imag} */,
  {32'hc4664e41, 32'h00000000} /* (27, 12, 0) {real, imag} */,
  {32'hc403ae97, 32'h432606b9} /* (27, 11, 31) {real, imag} */,
  {32'h439794eb, 32'h42565470} /* (27, 11, 30) {real, imag} */,
  {32'hc1b50110, 32'hc1afbbd0} /* (27, 11, 29) {real, imag} */,
  {32'hc1aea29c, 32'hc2fd3e0e} /* (27, 11, 28) {real, imag} */,
  {32'h4285f620, 32'hc29e75f7} /* (27, 11, 27) {real, imag} */,
  {32'h40266e50, 32'hc124d038} /* (27, 11, 26) {real, imag} */,
  {32'h424d847d, 32'hc27beef3} /* (27, 11, 25) {real, imag} */,
  {32'hc195a17c, 32'h419b6dfa} /* (27, 11, 24) {real, imag} */,
  {32'h415480da, 32'hc2922242} /* (27, 11, 23) {real, imag} */,
  {32'hc305a0b8, 32'h43196c01} /* (27, 11, 22) {real, imag} */,
  {32'h430098fb, 32'hc11da283} /* (27, 11, 21) {real, imag} */,
  {32'hc1e54792, 32'hc28142c7} /* (27, 11, 20) {real, imag} */,
  {32'h42345c0e, 32'hc1fb8657} /* (27, 11, 19) {real, imag} */,
  {32'h4226c280, 32'hc1284992} /* (27, 11, 18) {real, imag} */,
  {32'h41a5c8be, 32'h3fdb71e0} /* (27, 11, 17) {real, imag} */,
  {32'hc2313e66, 32'h00000000} /* (27, 11, 16) {real, imag} */,
  {32'h41a5c8be, 32'hbfdb71e0} /* (27, 11, 15) {real, imag} */,
  {32'h4226c280, 32'h41284992} /* (27, 11, 14) {real, imag} */,
  {32'h42345c0e, 32'h41fb8657} /* (27, 11, 13) {real, imag} */,
  {32'hc1e54792, 32'h428142c7} /* (27, 11, 12) {real, imag} */,
  {32'h430098fb, 32'h411da283} /* (27, 11, 11) {real, imag} */,
  {32'hc305a0b8, 32'hc3196c01} /* (27, 11, 10) {real, imag} */,
  {32'h415480da, 32'h42922242} /* (27, 11, 9) {real, imag} */,
  {32'hc195a17c, 32'hc19b6dfa} /* (27, 11, 8) {real, imag} */,
  {32'h424d847d, 32'h427beef3} /* (27, 11, 7) {real, imag} */,
  {32'h40266e50, 32'h4124d038} /* (27, 11, 6) {real, imag} */,
  {32'h4285f620, 32'h429e75f7} /* (27, 11, 5) {real, imag} */,
  {32'hc1aea29c, 32'h42fd3e0e} /* (27, 11, 4) {real, imag} */,
  {32'hc1b50110, 32'h41afbbd0} /* (27, 11, 3) {real, imag} */,
  {32'h439794eb, 32'hc2565470} /* (27, 11, 2) {real, imag} */,
  {32'hc403ae97, 32'hc32606b9} /* (27, 11, 1) {real, imag} */,
  {32'hc40d43ae, 32'h00000000} /* (27, 11, 0) {real, imag} */,
  {32'h43912615, 32'h431e40fc} /* (27, 10, 31) {real, imag} */,
  {32'hc388d130, 32'h432f9c69} /* (27, 10, 30) {real, imag} */,
  {32'hc2a55cc1, 32'h407a1b90} /* (27, 10, 29) {real, imag} */,
  {32'h43361509, 32'hc3a36414} /* (27, 10, 28) {real, imag} */,
  {32'h41c15d78, 32'h4302f1ab} /* (27, 10, 27) {real, imag} */,
  {32'h41a9e87c, 32'h41b42ea4} /* (27, 10, 26) {real, imag} */,
  {32'h4276d426, 32'hc295aa57} /* (27, 10, 25) {real, imag} */,
  {32'hc290d42d, 32'h42307aca} /* (27, 10, 24) {real, imag} */,
  {32'h41cc29c6, 32'h419dfe6c} /* (27, 10, 23) {real, imag} */,
  {32'h41e36bc8, 32'h4199d27c} /* (27, 10, 22) {real, imag} */,
  {32'h3f9f5a94, 32'h42a22b10} /* (27, 10, 21) {real, imag} */,
  {32'hc2bba63f, 32'hc1882d8c} /* (27, 10, 20) {real, imag} */,
  {32'h40966792, 32'hbf266040} /* (27, 10, 19) {real, imag} */,
  {32'hc24f295d, 32'h402fe640} /* (27, 10, 18) {real, imag} */,
  {32'hc115a378, 32'hc19b289c} /* (27, 10, 17) {real, imag} */,
  {32'h42aaf656, 32'h00000000} /* (27, 10, 16) {real, imag} */,
  {32'hc115a378, 32'h419b289c} /* (27, 10, 15) {real, imag} */,
  {32'hc24f295d, 32'hc02fe640} /* (27, 10, 14) {real, imag} */,
  {32'h40966792, 32'h3f266040} /* (27, 10, 13) {real, imag} */,
  {32'hc2bba63f, 32'h41882d8c} /* (27, 10, 12) {real, imag} */,
  {32'h3f9f5a94, 32'hc2a22b10} /* (27, 10, 11) {real, imag} */,
  {32'h41e36bc8, 32'hc199d27c} /* (27, 10, 10) {real, imag} */,
  {32'h41cc29c6, 32'hc19dfe6c} /* (27, 10, 9) {real, imag} */,
  {32'hc290d42d, 32'hc2307aca} /* (27, 10, 8) {real, imag} */,
  {32'h4276d426, 32'h4295aa57} /* (27, 10, 7) {real, imag} */,
  {32'h41a9e87c, 32'hc1b42ea4} /* (27, 10, 6) {real, imag} */,
  {32'h41c15d78, 32'hc302f1ab} /* (27, 10, 5) {real, imag} */,
  {32'h43361509, 32'h43a36414} /* (27, 10, 4) {real, imag} */,
  {32'hc2a55cc1, 32'hc07a1b90} /* (27, 10, 3) {real, imag} */,
  {32'hc388d130, 32'hc32f9c69} /* (27, 10, 2) {real, imag} */,
  {32'h43912615, 32'hc31e40fc} /* (27, 10, 1) {real, imag} */,
  {32'hc271fb7e, 32'h00000000} /* (27, 10, 0) {real, imag} */,
  {32'h443b520a, 32'h42ed7cb2} /* (27, 9, 31) {real, imag} */,
  {32'hc4044530, 32'h42f68f23} /* (27, 9, 30) {real, imag} */,
  {32'h4311542f, 32'hc27a2952} /* (27, 9, 29) {real, imag} */,
  {32'h433c35d9, 32'hc31e0422} /* (27, 9, 28) {real, imag} */,
  {32'hc340bba9, 32'h4277a3d6} /* (27, 9, 27) {real, imag} */,
  {32'h4254afa5, 32'h406f67e0} /* (27, 9, 26) {real, imag} */,
  {32'h4228839e, 32'hc1be3e9e} /* (27, 9, 25) {real, imag} */,
  {32'hc22be9ea, 32'h42afb762} /* (27, 9, 24) {real, imag} */,
  {32'h428685ad, 32'hc123f878} /* (27, 9, 23) {real, imag} */,
  {32'hc2444ea4, 32'hc245e57a} /* (27, 9, 22) {real, imag} */,
  {32'h422d6cb8, 32'h41d4a956} /* (27, 9, 21) {real, imag} */,
  {32'hc2052cba, 32'h418fe5ed} /* (27, 9, 20) {real, imag} */,
  {32'hc22c95c6, 32'h420a29fa} /* (27, 9, 19) {real, imag} */,
  {32'h42073c31, 32'h4215bfa0} /* (27, 9, 18) {real, imag} */,
  {32'hc261383b, 32'h40310a10} /* (27, 9, 17) {real, imag} */,
  {32'h42055efd, 32'h00000000} /* (27, 9, 16) {real, imag} */,
  {32'hc261383b, 32'hc0310a10} /* (27, 9, 15) {real, imag} */,
  {32'h42073c31, 32'hc215bfa0} /* (27, 9, 14) {real, imag} */,
  {32'hc22c95c6, 32'hc20a29fa} /* (27, 9, 13) {real, imag} */,
  {32'hc2052cba, 32'hc18fe5ed} /* (27, 9, 12) {real, imag} */,
  {32'h422d6cb8, 32'hc1d4a956} /* (27, 9, 11) {real, imag} */,
  {32'hc2444ea4, 32'h4245e57a} /* (27, 9, 10) {real, imag} */,
  {32'h428685ad, 32'h4123f878} /* (27, 9, 9) {real, imag} */,
  {32'hc22be9ea, 32'hc2afb762} /* (27, 9, 8) {real, imag} */,
  {32'h4228839e, 32'h41be3e9e} /* (27, 9, 7) {real, imag} */,
  {32'h4254afa5, 32'hc06f67e0} /* (27, 9, 6) {real, imag} */,
  {32'hc340bba9, 32'hc277a3d6} /* (27, 9, 5) {real, imag} */,
  {32'h433c35d9, 32'h431e0422} /* (27, 9, 4) {real, imag} */,
  {32'h4311542f, 32'h427a2952} /* (27, 9, 3) {real, imag} */,
  {32'hc4044530, 32'hc2f68f23} /* (27, 9, 2) {real, imag} */,
  {32'h443b520a, 32'hc2ed7cb2} /* (27, 9, 1) {real, imag} */,
  {32'h425ed294, 32'h00000000} /* (27, 9, 0) {real, imag} */,
  {32'h4463ca7f, 32'h4203bafb} /* (27, 8, 31) {real, imag} */,
  {32'hc42878df, 32'h438ee356} /* (27, 8, 30) {real, imag} */,
  {32'h4275ac39, 32'hc23c2c44} /* (27, 8, 29) {real, imag} */,
  {32'h4295a7e1, 32'hc347fff6} /* (27, 8, 28) {real, imag} */,
  {32'hc2fe36e3, 32'h42e697de} /* (27, 8, 27) {real, imag} */,
  {32'hc13cd664, 32'h4054e7c0} /* (27, 8, 26) {real, imag} */,
  {32'h41dda460, 32'hc2e34c94} /* (27, 8, 25) {real, imag} */,
  {32'hc2921118, 32'h432ef864} /* (27, 8, 24) {real, imag} */,
  {32'h42701ffb, 32'hc089ff88} /* (27, 8, 23) {real, imag} */,
  {32'h430b5356, 32'hc1797a64} /* (27, 8, 22) {real, imag} */,
  {32'h41e11e8e, 32'hc0b1fe10} /* (27, 8, 21) {real, imag} */,
  {32'h42233e60, 32'h42dc0099} /* (27, 8, 20) {real, imag} */,
  {32'h42b509c9, 32'hc2eeec8e} /* (27, 8, 19) {real, imag} */,
  {32'hc2b99ff9, 32'hc1e898d6} /* (27, 8, 18) {real, imag} */,
  {32'hc26b8f72, 32'h412b80cc} /* (27, 8, 17) {real, imag} */,
  {32'h416a68e6, 32'h00000000} /* (27, 8, 16) {real, imag} */,
  {32'hc26b8f72, 32'hc12b80cc} /* (27, 8, 15) {real, imag} */,
  {32'hc2b99ff9, 32'h41e898d6} /* (27, 8, 14) {real, imag} */,
  {32'h42b509c9, 32'h42eeec8e} /* (27, 8, 13) {real, imag} */,
  {32'h42233e60, 32'hc2dc0099} /* (27, 8, 12) {real, imag} */,
  {32'h41e11e8e, 32'h40b1fe10} /* (27, 8, 11) {real, imag} */,
  {32'h430b5356, 32'h41797a64} /* (27, 8, 10) {real, imag} */,
  {32'h42701ffb, 32'h4089ff88} /* (27, 8, 9) {real, imag} */,
  {32'hc2921118, 32'hc32ef864} /* (27, 8, 8) {real, imag} */,
  {32'h41dda460, 32'h42e34c94} /* (27, 8, 7) {real, imag} */,
  {32'hc13cd664, 32'hc054e7c0} /* (27, 8, 6) {real, imag} */,
  {32'hc2fe36e3, 32'hc2e697de} /* (27, 8, 5) {real, imag} */,
  {32'h4295a7e1, 32'h4347fff6} /* (27, 8, 4) {real, imag} */,
  {32'h4275ac39, 32'h423c2c44} /* (27, 8, 3) {real, imag} */,
  {32'hc42878df, 32'hc38ee356} /* (27, 8, 2) {real, imag} */,
  {32'h4463ca7f, 32'hc203bafb} /* (27, 8, 1) {real, imag} */,
  {32'hc24bb7ee, 32'h00000000} /* (27, 8, 0) {real, imag} */,
  {32'h445348ce, 32'h422e97c8} /* (27, 7, 31) {real, imag} */,
  {32'hc41bb884, 32'h43aec208} /* (27, 7, 30) {real, imag} */,
  {32'h415f7310, 32'h42c41a6e} /* (27, 7, 29) {real, imag} */,
  {32'h4253b3f4, 32'hc2c3aac2} /* (27, 7, 28) {real, imag} */,
  {32'hc242ef45, 32'h42a551f1} /* (27, 7, 27) {real, imag} */,
  {32'h41fe71ec, 32'hc1120fb0} /* (27, 7, 26) {real, imag} */,
  {32'h413c4bf8, 32'hc23ce63d} /* (27, 7, 25) {real, imag} */,
  {32'h4235cb14, 32'h41c6cdc3} /* (27, 7, 24) {real, imag} */,
  {32'hc22bac66, 32'h42a67210} /* (27, 7, 23) {real, imag} */,
  {32'hc2a13d80, 32'hc2b7551b} /* (27, 7, 22) {real, imag} */,
  {32'hc2787d62, 32'h414973d4} /* (27, 7, 21) {real, imag} */,
  {32'hc24a6d3e, 32'hc23d6346} /* (27, 7, 20) {real, imag} */,
  {32'h42384504, 32'h41d4648e} /* (27, 7, 19) {real, imag} */,
  {32'h42d87db4, 32'hc13e9c78} /* (27, 7, 18) {real, imag} */,
  {32'hc1a27700, 32'h411de454} /* (27, 7, 17) {real, imag} */,
  {32'hc2158052, 32'h00000000} /* (27, 7, 16) {real, imag} */,
  {32'hc1a27700, 32'hc11de454} /* (27, 7, 15) {real, imag} */,
  {32'h42d87db4, 32'h413e9c78} /* (27, 7, 14) {real, imag} */,
  {32'h42384504, 32'hc1d4648e} /* (27, 7, 13) {real, imag} */,
  {32'hc24a6d3e, 32'h423d6346} /* (27, 7, 12) {real, imag} */,
  {32'hc2787d62, 32'hc14973d4} /* (27, 7, 11) {real, imag} */,
  {32'hc2a13d80, 32'h42b7551b} /* (27, 7, 10) {real, imag} */,
  {32'hc22bac66, 32'hc2a67210} /* (27, 7, 9) {real, imag} */,
  {32'h4235cb14, 32'hc1c6cdc3} /* (27, 7, 8) {real, imag} */,
  {32'h413c4bf8, 32'h423ce63d} /* (27, 7, 7) {real, imag} */,
  {32'h41fe71ec, 32'h41120fb0} /* (27, 7, 6) {real, imag} */,
  {32'hc242ef45, 32'hc2a551f1} /* (27, 7, 5) {real, imag} */,
  {32'h4253b3f4, 32'h42c3aac2} /* (27, 7, 4) {real, imag} */,
  {32'h415f7310, 32'hc2c41a6e} /* (27, 7, 3) {real, imag} */,
  {32'hc41bb884, 32'hc3aec208} /* (27, 7, 2) {real, imag} */,
  {32'h445348ce, 32'hc22e97c8} /* (27, 7, 1) {real, imag} */,
  {32'hc2851d22, 32'h00000000} /* (27, 7, 0) {real, imag} */,
  {32'h442859eb, 32'h41957d80} /* (27, 6, 31) {real, imag} */,
  {32'hc40a8320, 32'h43d162c2} /* (27, 6, 30) {real, imag} */,
  {32'hbfb8b0f0, 32'h40a96860} /* (27, 6, 29) {real, imag} */,
  {32'h43041c7c, 32'h4244de3e} /* (27, 6, 28) {real, imag} */,
  {32'hc30ade04, 32'h42dc0c10} /* (27, 6, 27) {real, imag} */,
  {32'h4354c4ca, 32'hc29df57d} /* (27, 6, 26) {real, imag} */,
  {32'hc2575d90, 32'h417c2056} /* (27, 6, 25) {real, imag} */,
  {32'hc1483939, 32'h43153372} /* (27, 6, 24) {real, imag} */,
  {32'hc1c34f96, 32'h425a09b8} /* (27, 6, 23) {real, imag} */,
  {32'hc2087c17, 32'hc100555e} /* (27, 6, 22) {real, imag} */,
  {32'hc1eb949f, 32'h42bd1762} /* (27, 6, 21) {real, imag} */,
  {32'hc289fcf4, 32'h42483ef4} /* (27, 6, 20) {real, imag} */,
  {32'h40973810, 32'hc2b55e77} /* (27, 6, 19) {real, imag} */,
  {32'h4219022b, 32'h42913b88} /* (27, 6, 18) {real, imag} */,
  {32'hc246043f, 32'hc187e8f8} /* (27, 6, 17) {real, imag} */,
  {32'hc287b651, 32'h00000000} /* (27, 6, 16) {real, imag} */,
  {32'hc246043f, 32'h4187e8f8} /* (27, 6, 15) {real, imag} */,
  {32'h4219022b, 32'hc2913b88} /* (27, 6, 14) {real, imag} */,
  {32'h40973810, 32'h42b55e77} /* (27, 6, 13) {real, imag} */,
  {32'hc289fcf4, 32'hc2483ef4} /* (27, 6, 12) {real, imag} */,
  {32'hc1eb949f, 32'hc2bd1762} /* (27, 6, 11) {real, imag} */,
  {32'hc2087c17, 32'h4100555e} /* (27, 6, 10) {real, imag} */,
  {32'hc1c34f96, 32'hc25a09b8} /* (27, 6, 9) {real, imag} */,
  {32'hc1483939, 32'hc3153372} /* (27, 6, 8) {real, imag} */,
  {32'hc2575d90, 32'hc17c2056} /* (27, 6, 7) {real, imag} */,
  {32'h4354c4ca, 32'h429df57d} /* (27, 6, 6) {real, imag} */,
  {32'hc30ade04, 32'hc2dc0c10} /* (27, 6, 5) {real, imag} */,
  {32'h43041c7c, 32'hc244de3e} /* (27, 6, 4) {real, imag} */,
  {32'hbfb8b0f0, 32'hc0a96860} /* (27, 6, 3) {real, imag} */,
  {32'hc40a8320, 32'hc3d162c2} /* (27, 6, 2) {real, imag} */,
  {32'h442859eb, 32'hc1957d80} /* (27, 6, 1) {real, imag} */,
  {32'h42360520, 32'h00000000} /* (27, 6, 0) {real, imag} */,
  {32'h43bd6982, 32'hc399f415} /* (27, 5, 31) {real, imag} */,
  {32'hc38596b9, 32'h43e18222} /* (27, 5, 30) {real, imag} */,
  {32'h41826b70, 32'hc1930627} /* (27, 5, 29) {real, imag} */,
  {32'hc1954aa2, 32'h42ecbd56} /* (27, 5, 28) {real, imag} */,
  {32'hc2cf0fd0, 32'h421956ce} /* (27, 5, 27) {real, imag} */,
  {32'h4288056e, 32'hc291827f} /* (27, 5, 26) {real, imag} */,
  {32'hc2d5ec3e, 32'h4189ff89} /* (27, 5, 25) {real, imag} */,
  {32'hc1c27db3, 32'h4308cb82} /* (27, 5, 24) {real, imag} */,
  {32'hc0e6a9fe, 32'h413f79a8} /* (27, 5, 23) {real, imag} */,
  {32'h426d92a1, 32'hc29e8cd0} /* (27, 5, 22) {real, imag} */,
  {32'hc1c62840, 32'h41fd9656} /* (27, 5, 21) {real, imag} */,
  {32'hc2400858, 32'h4177126c} /* (27, 5, 20) {real, imag} */,
  {32'h42b8f228, 32'h41a73b30} /* (27, 5, 19) {real, imag} */,
  {32'hc15fe3f7, 32'hc2282f48} /* (27, 5, 18) {real, imag} */,
  {32'h4205df32, 32'h42102ff9} /* (27, 5, 17) {real, imag} */,
  {32'h419aef7b, 32'h00000000} /* (27, 5, 16) {real, imag} */,
  {32'h4205df32, 32'hc2102ff9} /* (27, 5, 15) {real, imag} */,
  {32'hc15fe3f7, 32'h42282f48} /* (27, 5, 14) {real, imag} */,
  {32'h42b8f228, 32'hc1a73b30} /* (27, 5, 13) {real, imag} */,
  {32'hc2400858, 32'hc177126c} /* (27, 5, 12) {real, imag} */,
  {32'hc1c62840, 32'hc1fd9656} /* (27, 5, 11) {real, imag} */,
  {32'h426d92a1, 32'h429e8cd0} /* (27, 5, 10) {real, imag} */,
  {32'hc0e6a9fe, 32'hc13f79a8} /* (27, 5, 9) {real, imag} */,
  {32'hc1c27db3, 32'hc308cb82} /* (27, 5, 8) {real, imag} */,
  {32'hc2d5ec3e, 32'hc189ff89} /* (27, 5, 7) {real, imag} */,
  {32'h4288056e, 32'h4291827f} /* (27, 5, 6) {real, imag} */,
  {32'hc2cf0fd0, 32'hc21956ce} /* (27, 5, 5) {real, imag} */,
  {32'hc1954aa2, 32'hc2ecbd56} /* (27, 5, 4) {real, imag} */,
  {32'h41826b70, 32'h41930627} /* (27, 5, 3) {real, imag} */,
  {32'hc38596b9, 32'hc3e18222} /* (27, 5, 2) {real, imag} */,
  {32'h43bd6982, 32'h4399f415} /* (27, 5, 1) {real, imag} */,
  {32'hc1a60960, 32'h00000000} /* (27, 5, 0) {real, imag} */,
  {32'h428e1dd0, 32'hc3b6797f} /* (27, 4, 31) {real, imag} */,
  {32'h43171454, 32'h442dff03} /* (27, 4, 30) {real, imag} */,
  {32'hc2ddbbe0, 32'hc0c1da70} /* (27, 4, 29) {real, imag} */,
  {32'hc2fec6a6, 32'h420485a8} /* (27, 4, 28) {real, imag} */,
  {32'hc3848578, 32'hc2540b79} /* (27, 4, 27) {real, imag} */,
  {32'h42805696, 32'h42262331} /* (27, 4, 26) {real, imag} */,
  {32'h41caafb8, 32'hc13a4a38} /* (27, 4, 25) {real, imag} */,
  {32'h42e1bb0d, 32'h41b32c5c} /* (27, 4, 24) {real, imag} */,
  {32'hc2938c6d, 32'hc21dc577} /* (27, 4, 23) {real, imag} */,
  {32'hc20257c6, 32'h413db4fa} /* (27, 4, 22) {real, imag} */,
  {32'hbf1d5440, 32'hc2361dea} /* (27, 4, 21) {real, imag} */,
  {32'hc24f183a, 32'h4045c720} /* (27, 4, 20) {real, imag} */,
  {32'h4282d7fe, 32'hc0a61870} /* (27, 4, 19) {real, imag} */,
  {32'h42747cda, 32'h4200bb14} /* (27, 4, 18) {real, imag} */,
  {32'hc25a6872, 32'h42ad6c10} /* (27, 4, 17) {real, imag} */,
  {32'h40f59584, 32'h00000000} /* (27, 4, 16) {real, imag} */,
  {32'hc25a6872, 32'hc2ad6c10} /* (27, 4, 15) {real, imag} */,
  {32'h42747cda, 32'hc200bb14} /* (27, 4, 14) {real, imag} */,
  {32'h4282d7fe, 32'h40a61870} /* (27, 4, 13) {real, imag} */,
  {32'hc24f183a, 32'hc045c720} /* (27, 4, 12) {real, imag} */,
  {32'hbf1d5440, 32'h42361dea} /* (27, 4, 11) {real, imag} */,
  {32'hc20257c6, 32'hc13db4fa} /* (27, 4, 10) {real, imag} */,
  {32'hc2938c6d, 32'h421dc577} /* (27, 4, 9) {real, imag} */,
  {32'h42e1bb0d, 32'hc1b32c5c} /* (27, 4, 8) {real, imag} */,
  {32'h41caafb8, 32'h413a4a38} /* (27, 4, 7) {real, imag} */,
  {32'h42805696, 32'hc2262331} /* (27, 4, 6) {real, imag} */,
  {32'hc3848578, 32'h42540b79} /* (27, 4, 5) {real, imag} */,
  {32'hc2fec6a6, 32'hc20485a8} /* (27, 4, 4) {real, imag} */,
  {32'hc2ddbbe0, 32'h40c1da70} /* (27, 4, 3) {real, imag} */,
  {32'h43171454, 32'hc42dff03} /* (27, 4, 2) {real, imag} */,
  {32'h428e1dd0, 32'h43b6797f} /* (27, 4, 1) {real, imag} */,
  {32'hc31be3c8, 32'h00000000} /* (27, 4, 0) {real, imag} */,
  {32'hc1ecb570, 32'hc4111ea5} /* (27, 3, 31) {real, imag} */,
  {32'h43943e09, 32'h441664c2} /* (27, 3, 30) {real, imag} */,
  {32'hc2a30f74, 32'hc2c73a56} /* (27, 3, 29) {real, imag} */,
  {32'hc2d4971e, 32'h42b2ee87} /* (27, 3, 28) {real, imag} */,
  {32'hc319b458, 32'h423bb877} /* (27, 3, 27) {real, imag} */,
  {32'hc21e7b96, 32'h41a0111c} /* (27, 3, 26) {real, imag} */,
  {32'h40420f30, 32'h42424dee} /* (27, 3, 25) {real, imag} */,
  {32'h416d41a8, 32'h4242a7eb} /* (27, 3, 24) {real, imag} */,
  {32'hc1a8ed6d, 32'h41aea8da} /* (27, 3, 23) {real, imag} */,
  {32'hc2b906fb, 32'h424d481a} /* (27, 3, 22) {real, imag} */,
  {32'h417c4b34, 32'hc1f06082} /* (27, 3, 21) {real, imag} */,
  {32'h4205f899, 32'h428721bf} /* (27, 3, 20) {real, imag} */,
  {32'h41c32bea, 32'hc2090726} /* (27, 3, 19) {real, imag} */,
  {32'h429a9f06, 32'h429b3a12} /* (27, 3, 18) {real, imag} */,
  {32'hc0c306e8, 32'hc277bda7} /* (27, 3, 17) {real, imag} */,
  {32'h42003a29, 32'h00000000} /* (27, 3, 16) {real, imag} */,
  {32'hc0c306e8, 32'h4277bda7} /* (27, 3, 15) {real, imag} */,
  {32'h429a9f06, 32'hc29b3a12} /* (27, 3, 14) {real, imag} */,
  {32'h41c32bea, 32'h42090726} /* (27, 3, 13) {real, imag} */,
  {32'h4205f899, 32'hc28721bf} /* (27, 3, 12) {real, imag} */,
  {32'h417c4b34, 32'h41f06082} /* (27, 3, 11) {real, imag} */,
  {32'hc2b906fb, 32'hc24d481a} /* (27, 3, 10) {real, imag} */,
  {32'hc1a8ed6d, 32'hc1aea8da} /* (27, 3, 9) {real, imag} */,
  {32'h416d41a8, 32'hc242a7eb} /* (27, 3, 8) {real, imag} */,
  {32'h40420f30, 32'hc2424dee} /* (27, 3, 7) {real, imag} */,
  {32'hc21e7b96, 32'hc1a0111c} /* (27, 3, 6) {real, imag} */,
  {32'hc319b458, 32'hc23bb877} /* (27, 3, 5) {real, imag} */,
  {32'hc2d4971e, 32'hc2b2ee87} /* (27, 3, 4) {real, imag} */,
  {32'hc2a30f74, 32'h42c73a56} /* (27, 3, 3) {real, imag} */,
  {32'h43943e09, 32'hc41664c2} /* (27, 3, 2) {real, imag} */,
  {32'hc1ecb570, 32'h44111ea5} /* (27, 3, 1) {real, imag} */,
  {32'hc29abbc4, 32'h00000000} /* (27, 3, 0) {real, imag} */,
  {32'hc2f9eaec, 32'hc43e19e0} /* (27, 2, 31) {real, imag} */,
  {32'h43bae610, 32'h442669c1} /* (27, 2, 30) {real, imag} */,
  {32'hc1c70c28, 32'hc15da488} /* (27, 2, 29) {real, imag} */,
  {32'hc28924ba, 32'h4308cd05} /* (27, 2, 28) {real, imag} */,
  {32'hc2925bd9, 32'h428ce3be} /* (27, 2, 27) {real, imag} */,
  {32'hc20c14de, 32'h42aac6be} /* (27, 2, 26) {real, imag} */,
  {32'hc2dcf206, 32'hc1b590ff} /* (27, 2, 25) {real, imag} */,
  {32'h428d3ae2, 32'h42838e00} /* (27, 2, 24) {real, imag} */,
  {32'hc2931d5f, 32'hc23e0a0a} /* (27, 2, 23) {real, imag} */,
  {32'hc1759622, 32'h42e781f4} /* (27, 2, 22) {real, imag} */,
  {32'hc2c4c62e, 32'h411046ce} /* (27, 2, 21) {real, imag} */,
  {32'h42a2bb59, 32'h4219a95a} /* (27, 2, 20) {real, imag} */,
  {32'hc23d8530, 32'hc2b49d66} /* (27, 2, 19) {real, imag} */,
  {32'h421f8482, 32'h42daa3de} /* (27, 2, 18) {real, imag} */,
  {32'h424b1db8, 32'h41d08bd3} /* (27, 2, 17) {real, imag} */,
  {32'hc1c00ec0, 32'h00000000} /* (27, 2, 16) {real, imag} */,
  {32'h424b1db8, 32'hc1d08bd3} /* (27, 2, 15) {real, imag} */,
  {32'h421f8482, 32'hc2daa3de} /* (27, 2, 14) {real, imag} */,
  {32'hc23d8530, 32'h42b49d66} /* (27, 2, 13) {real, imag} */,
  {32'h42a2bb59, 32'hc219a95a} /* (27, 2, 12) {real, imag} */,
  {32'hc2c4c62e, 32'hc11046ce} /* (27, 2, 11) {real, imag} */,
  {32'hc1759622, 32'hc2e781f4} /* (27, 2, 10) {real, imag} */,
  {32'hc2931d5f, 32'h423e0a0a} /* (27, 2, 9) {real, imag} */,
  {32'h428d3ae2, 32'hc2838e00} /* (27, 2, 8) {real, imag} */,
  {32'hc2dcf206, 32'h41b590ff} /* (27, 2, 7) {real, imag} */,
  {32'hc20c14de, 32'hc2aac6be} /* (27, 2, 6) {real, imag} */,
  {32'hc2925bd9, 32'hc28ce3be} /* (27, 2, 5) {real, imag} */,
  {32'hc28924ba, 32'hc308cd05} /* (27, 2, 4) {real, imag} */,
  {32'hc1c70c28, 32'h415da488} /* (27, 2, 3) {real, imag} */,
  {32'h43bae610, 32'hc42669c1} /* (27, 2, 2) {real, imag} */,
  {32'hc2f9eaec, 32'h443e19e0} /* (27, 2, 1) {real, imag} */,
  {32'hc370427a, 32'h00000000} /* (27, 2, 0) {real, imag} */,
  {32'hc2e45e12, 32'hc456e2b8} /* (27, 1, 31) {real, imag} */,
  {32'h43e5d5ea, 32'h442b7416} /* (27, 1, 30) {real, imag} */,
  {32'hc10b85e8, 32'hc140dcde} /* (27, 1, 29) {real, imag} */,
  {32'h41ea2a34, 32'h42dcfacc} /* (27, 1, 28) {real, imag} */,
  {32'hc2d5b77d, 32'hc2e1e79c} /* (27, 1, 27) {real, imag} */,
  {32'h421f323a, 32'h4288ba94} /* (27, 1, 26) {real, imag} */,
  {32'hc21a48d2, 32'hc19d62ff} /* (27, 1, 25) {real, imag} */,
  {32'hc2b7bf3e, 32'h422b4dac} /* (27, 1, 24) {real, imag} */,
  {32'hc16c2922, 32'h3e6ac700} /* (27, 1, 23) {real, imag} */,
  {32'h42436009, 32'h420f9a78} /* (27, 1, 22) {real, imag} */,
  {32'hc3382c62, 32'h42ace78c} /* (27, 1, 21) {real, imag} */,
  {32'h423ba695, 32'h427a37b8} /* (27, 1, 20) {real, imag} */,
  {32'h426f1d80, 32'hc00fec2c} /* (27, 1, 19) {real, imag} */,
  {32'h42aadf5e, 32'hc14a831a} /* (27, 1, 18) {real, imag} */,
  {32'hc16d72d8, 32'hc23ea032} /* (27, 1, 17) {real, imag} */,
  {32'hc26c3d1c, 32'h00000000} /* (27, 1, 16) {real, imag} */,
  {32'hc16d72d8, 32'h423ea032} /* (27, 1, 15) {real, imag} */,
  {32'h42aadf5e, 32'h414a831a} /* (27, 1, 14) {real, imag} */,
  {32'h426f1d80, 32'h400fec2c} /* (27, 1, 13) {real, imag} */,
  {32'h423ba695, 32'hc27a37b8} /* (27, 1, 12) {real, imag} */,
  {32'hc3382c62, 32'hc2ace78c} /* (27, 1, 11) {real, imag} */,
  {32'h42436009, 32'hc20f9a78} /* (27, 1, 10) {real, imag} */,
  {32'hc16c2922, 32'hbe6ac700} /* (27, 1, 9) {real, imag} */,
  {32'hc2b7bf3e, 32'hc22b4dac} /* (27, 1, 8) {real, imag} */,
  {32'hc21a48d2, 32'h419d62ff} /* (27, 1, 7) {real, imag} */,
  {32'h421f323a, 32'hc288ba94} /* (27, 1, 6) {real, imag} */,
  {32'hc2d5b77d, 32'h42e1e79c} /* (27, 1, 5) {real, imag} */,
  {32'h41ea2a34, 32'hc2dcfacc} /* (27, 1, 4) {real, imag} */,
  {32'hc10b85e8, 32'h4140dcde} /* (27, 1, 3) {real, imag} */,
  {32'h43e5d5ea, 32'hc42b7416} /* (27, 1, 2) {real, imag} */,
  {32'hc2e45e12, 32'h4456e2b8} /* (27, 1, 1) {real, imag} */,
  {32'hc3988256, 32'h00000000} /* (27, 1, 0) {real, imag} */,
  {32'hc35e3664, 32'hc3c00c76} /* (27, 0, 31) {real, imag} */,
  {32'h429a2608, 32'h43eee51a} /* (27, 0, 30) {real, imag} */,
  {32'h40dfa408, 32'hc214ea6e} /* (27, 0, 29) {real, imag} */,
  {32'hc0a32db0, 32'h431bd077} /* (27, 0, 28) {real, imag} */,
  {32'hc3002aae, 32'hc2a701bc} /* (27, 0, 27) {real, imag} */,
  {32'hc28bd4e2, 32'h411c634b} /* (27, 0, 26) {real, imag} */,
  {32'h4297f8e0, 32'hc273b1cd} /* (27, 0, 25) {real, imag} */,
  {32'hc2a3db55, 32'h3febe300} /* (27, 0, 24) {real, imag} */,
  {32'h4246ddd5, 32'h42147a34} /* (27, 0, 23) {real, imag} */,
  {32'h41202ea8, 32'hc2018563} /* (27, 0, 22) {real, imag} */,
  {32'h40a86f44, 32'h42229fc6} /* (27, 0, 21) {real, imag} */,
  {32'h41b87dbb, 32'h418ac761} /* (27, 0, 20) {real, imag} */,
  {32'h40f19d7d, 32'hc10faf24} /* (27, 0, 19) {real, imag} */,
  {32'h41b037c5, 32'hc18f4794} /* (27, 0, 18) {real, imag} */,
  {32'hc1dd4e26, 32'h42528134} /* (27, 0, 17) {real, imag} */,
  {32'hc134c1eb, 32'h00000000} /* (27, 0, 16) {real, imag} */,
  {32'hc1dd4e26, 32'hc2528134} /* (27, 0, 15) {real, imag} */,
  {32'h41b037c5, 32'h418f4794} /* (27, 0, 14) {real, imag} */,
  {32'h40f19d7d, 32'h410faf24} /* (27, 0, 13) {real, imag} */,
  {32'h41b87dbb, 32'hc18ac761} /* (27, 0, 12) {real, imag} */,
  {32'h40a86f44, 32'hc2229fc6} /* (27, 0, 11) {real, imag} */,
  {32'h41202ea8, 32'h42018563} /* (27, 0, 10) {real, imag} */,
  {32'h4246ddd5, 32'hc2147a34} /* (27, 0, 9) {real, imag} */,
  {32'hc2a3db55, 32'hbfebe300} /* (27, 0, 8) {real, imag} */,
  {32'h4297f8e0, 32'h4273b1cd} /* (27, 0, 7) {real, imag} */,
  {32'hc28bd4e2, 32'hc11c634b} /* (27, 0, 6) {real, imag} */,
  {32'hc3002aae, 32'h42a701bc} /* (27, 0, 5) {real, imag} */,
  {32'hc0a32db0, 32'hc31bd077} /* (27, 0, 4) {real, imag} */,
  {32'h40dfa408, 32'h4214ea6e} /* (27, 0, 3) {real, imag} */,
  {32'h429a2608, 32'hc3eee51a} /* (27, 0, 2) {real, imag} */,
  {32'hc35e3664, 32'h43c00c76} /* (27, 0, 1) {real, imag} */,
  {32'hc41b3cfa, 32'h00000000} /* (27, 0, 0) {real, imag} */,
  {32'hc452a408, 32'h440ba03f} /* (26, 31, 31) {real, imag} */,
  {32'h42981b33, 32'h42c49ad2} /* (26, 31, 30) {real, imag} */,
  {32'hc2a1b7f2, 32'h41f3116a} /* (26, 31, 29) {real, imag} */,
  {32'h4253bfee, 32'h43072451} /* (26, 31, 28) {real, imag} */,
  {32'h422832a8, 32'hc21fb3ea} /* (26, 31, 27) {real, imag} */,
  {32'h42978668, 32'h42ca170c} /* (26, 31, 26) {real, imag} */,
  {32'h424b0762, 32'h419f162e} /* (26, 31, 25) {real, imag} */,
  {32'hc128c4c8, 32'hc0448d20} /* (26, 31, 24) {real, imag} */,
  {32'h41bfafa2, 32'h41a95af7} /* (26, 31, 23) {real, imag} */,
  {32'hc08f5fc4, 32'hc2b28dc6} /* (26, 31, 22) {real, imag} */,
  {32'h4187182c, 32'h426b9498} /* (26, 31, 21) {real, imag} */,
  {32'h42ba617b, 32'hc1f9f778} /* (26, 31, 20) {real, imag} */,
  {32'h428bcc14, 32'hc28729de} /* (26, 31, 19) {real, imag} */,
  {32'hbf9e61b0, 32'h4283d30e} /* (26, 31, 18) {real, imag} */,
  {32'h41469201, 32'h409d3844} /* (26, 31, 17) {real, imag} */,
  {32'hc28a5019, 32'h00000000} /* (26, 31, 16) {real, imag} */,
  {32'h41469201, 32'hc09d3844} /* (26, 31, 15) {real, imag} */,
  {32'hbf9e61b0, 32'hc283d30e} /* (26, 31, 14) {real, imag} */,
  {32'h428bcc14, 32'h428729de} /* (26, 31, 13) {real, imag} */,
  {32'h42ba617b, 32'h41f9f778} /* (26, 31, 12) {real, imag} */,
  {32'h4187182c, 32'hc26b9498} /* (26, 31, 11) {real, imag} */,
  {32'hc08f5fc4, 32'h42b28dc6} /* (26, 31, 10) {real, imag} */,
  {32'h41bfafa2, 32'hc1a95af7} /* (26, 31, 9) {real, imag} */,
  {32'hc128c4c8, 32'h40448d20} /* (26, 31, 8) {real, imag} */,
  {32'h424b0762, 32'hc19f162e} /* (26, 31, 7) {real, imag} */,
  {32'h42978668, 32'hc2ca170c} /* (26, 31, 6) {real, imag} */,
  {32'h422832a8, 32'h421fb3ea} /* (26, 31, 5) {real, imag} */,
  {32'h4253bfee, 32'hc3072451} /* (26, 31, 4) {real, imag} */,
  {32'hc2a1b7f2, 32'hc1f3116a} /* (26, 31, 3) {real, imag} */,
  {32'h42981b33, 32'hc2c49ad2} /* (26, 31, 2) {real, imag} */,
  {32'hc452a408, 32'hc40ba03f} /* (26, 31, 1) {real, imag} */,
  {32'hc4e70ef1, 32'h00000000} /* (26, 31, 0) {real, imag} */,
  {32'hc44a1c0b, 32'h43f3b043} /* (26, 30, 31) {real, imag} */,
  {32'h40c77e90, 32'h431ecf14} /* (26, 30, 30) {real, imag} */,
  {32'hc2f0fc6c, 32'hc17b8ef6} /* (26, 30, 29) {real, imag} */,
  {32'hc2b4754c, 32'h411715c9} /* (26, 30, 28) {real, imag} */,
  {32'hc1010c60, 32'hc2bd318f} /* (26, 30, 27) {real, imag} */,
  {32'h42a0a660, 32'h4211b2a6} /* (26, 30, 26) {real, imag} */,
  {32'h42505db4, 32'h427285ce} /* (26, 30, 25) {real, imag} */,
  {32'hc28fcb72, 32'hc2a83490} /* (26, 30, 24) {real, imag} */,
  {32'hc1e11a3e, 32'hc223867a} /* (26, 30, 23) {real, imag} */,
  {32'h3f0b1b90, 32'hc1877898} /* (26, 30, 22) {real, imag} */,
  {32'h4130ef74, 32'h42f9c3ee} /* (26, 30, 21) {real, imag} */,
  {32'h410ea896, 32'hc29d5c26} /* (26, 30, 20) {real, imag} */,
  {32'h419f5c5d, 32'h41f185e9} /* (26, 30, 19) {real, imag} */,
  {32'h420c60df, 32'hc2737058} /* (26, 30, 18) {real, imag} */,
  {32'hc1ca1767, 32'hc2852262} /* (26, 30, 17) {real, imag} */,
  {32'h428d9922, 32'h00000000} /* (26, 30, 16) {real, imag} */,
  {32'hc1ca1767, 32'h42852262} /* (26, 30, 15) {real, imag} */,
  {32'h420c60df, 32'h42737058} /* (26, 30, 14) {real, imag} */,
  {32'h419f5c5d, 32'hc1f185e9} /* (26, 30, 13) {real, imag} */,
  {32'h410ea896, 32'h429d5c26} /* (26, 30, 12) {real, imag} */,
  {32'h4130ef74, 32'hc2f9c3ee} /* (26, 30, 11) {real, imag} */,
  {32'h3f0b1b90, 32'h41877898} /* (26, 30, 10) {real, imag} */,
  {32'hc1e11a3e, 32'h4223867a} /* (26, 30, 9) {real, imag} */,
  {32'hc28fcb72, 32'h42a83490} /* (26, 30, 8) {real, imag} */,
  {32'h42505db4, 32'hc27285ce} /* (26, 30, 7) {real, imag} */,
  {32'h42a0a660, 32'hc211b2a6} /* (26, 30, 6) {real, imag} */,
  {32'hc1010c60, 32'h42bd318f} /* (26, 30, 5) {real, imag} */,
  {32'hc2b4754c, 32'hc11715c9} /* (26, 30, 4) {real, imag} */,
  {32'hc2f0fc6c, 32'h417b8ef6} /* (26, 30, 3) {real, imag} */,
  {32'h40c77e90, 32'hc31ecf14} /* (26, 30, 2) {real, imag} */,
  {32'hc44a1c0b, 32'hc3f3b043} /* (26, 30, 1) {real, imag} */,
  {32'hc4d7665c, 32'h00000000} /* (26, 30, 0) {real, imag} */,
  {32'hc43132f3, 32'h440751f9} /* (26, 29, 31) {real, imag} */,
  {32'hc24f7fc4, 32'h43235a1a} /* (26, 29, 30) {real, imag} */,
  {32'hc246a39e, 32'hc31530b4} /* (26, 29, 29) {real, imag} */,
  {32'hc18feea2, 32'hc27bc4b3} /* (26, 29, 28) {real, imag} */,
  {32'hc226e4af, 32'hc219c4b3} /* (26, 29, 27) {real, imag} */,
  {32'h40d30fe8, 32'hc3408204} /* (26, 29, 26) {real, imag} */,
  {32'h432e2964, 32'h40b8a67c} /* (26, 29, 25) {real, imag} */,
  {32'hc212c30d, 32'hc24cffa8} /* (26, 29, 24) {real, imag} */,
  {32'hc327881d, 32'hc2f78245} /* (26, 29, 23) {real, imag} */,
  {32'hc2677c6f, 32'hc203a888} /* (26, 29, 22) {real, imag} */,
  {32'hc233bfc4, 32'hc1154690} /* (26, 29, 21) {real, imag} */,
  {32'hc23dc636, 32'hc1bfdefb} /* (26, 29, 20) {real, imag} */,
  {32'h41cab38a, 32'hc1201268} /* (26, 29, 19) {real, imag} */,
  {32'h419540a0, 32'h42247a21} /* (26, 29, 18) {real, imag} */,
  {32'h41bf0c3a, 32'h41067d88} /* (26, 29, 17) {real, imag} */,
  {32'h41213c14, 32'h00000000} /* (26, 29, 16) {real, imag} */,
  {32'h41bf0c3a, 32'hc1067d88} /* (26, 29, 15) {real, imag} */,
  {32'h419540a0, 32'hc2247a21} /* (26, 29, 14) {real, imag} */,
  {32'h41cab38a, 32'h41201268} /* (26, 29, 13) {real, imag} */,
  {32'hc23dc636, 32'h41bfdefb} /* (26, 29, 12) {real, imag} */,
  {32'hc233bfc4, 32'h41154690} /* (26, 29, 11) {real, imag} */,
  {32'hc2677c6f, 32'h4203a888} /* (26, 29, 10) {real, imag} */,
  {32'hc327881d, 32'h42f78245} /* (26, 29, 9) {real, imag} */,
  {32'hc212c30d, 32'h424cffa8} /* (26, 29, 8) {real, imag} */,
  {32'h432e2964, 32'hc0b8a67c} /* (26, 29, 7) {real, imag} */,
  {32'h40d30fe8, 32'h43408204} /* (26, 29, 6) {real, imag} */,
  {32'hc226e4af, 32'h4219c4b3} /* (26, 29, 5) {real, imag} */,
  {32'hc18feea2, 32'h427bc4b3} /* (26, 29, 4) {real, imag} */,
  {32'hc246a39e, 32'h431530b4} /* (26, 29, 3) {real, imag} */,
  {32'hc24f7fc4, 32'hc3235a1a} /* (26, 29, 2) {real, imag} */,
  {32'hc43132f3, 32'hc40751f9} /* (26, 29, 1) {real, imag} */,
  {32'hc4e32cdb, 32'h00000000} /* (26, 29, 0) {real, imag} */,
  {32'hc425bc40, 32'h440c1cdf} /* (26, 28, 31) {real, imag} */,
  {32'hc2d9a4bf, 32'h4307b51e} /* (26, 28, 30) {real, imag} */,
  {32'h42a140f4, 32'hc3352b96} /* (26, 28, 29) {real, imag} */,
  {32'h42699df1, 32'hc1a6ceb6} /* (26, 28, 28) {real, imag} */,
  {32'h423fdaf3, 32'hc2851dee} /* (26, 28, 27) {real, imag} */,
  {32'h42b8c25b, 32'h4334c8e8} /* (26, 28, 26) {real, imag} */,
  {32'h431125f0, 32'hc2005a54} /* (26, 28, 25) {real, imag} */,
  {32'h3f94b580, 32'h4180f63c} /* (26, 28, 24) {real, imag} */,
  {32'hc1d56f90, 32'hc30cd4a8} /* (26, 28, 23) {real, imag} */,
  {32'hc3178ae4, 32'h423a531a} /* (26, 28, 22) {real, imag} */,
  {32'h4209a594, 32'h408a5638} /* (26, 28, 21) {real, imag} */,
  {32'h413d904e, 32'h43073983} /* (26, 28, 20) {real, imag} */,
  {32'hc1a7d5b4, 32'hc27b4d69} /* (26, 28, 19) {real, imag} */,
  {32'h41ebcfd5, 32'h42870926} /* (26, 28, 18) {real, imag} */,
  {32'h423a906f, 32'hc2651f14} /* (26, 28, 17) {real, imag} */,
  {32'h42ba4bc4, 32'h00000000} /* (26, 28, 16) {real, imag} */,
  {32'h423a906f, 32'h42651f14} /* (26, 28, 15) {real, imag} */,
  {32'h41ebcfd5, 32'hc2870926} /* (26, 28, 14) {real, imag} */,
  {32'hc1a7d5b4, 32'h427b4d69} /* (26, 28, 13) {real, imag} */,
  {32'h413d904e, 32'hc3073983} /* (26, 28, 12) {real, imag} */,
  {32'h4209a594, 32'hc08a5638} /* (26, 28, 11) {real, imag} */,
  {32'hc3178ae4, 32'hc23a531a} /* (26, 28, 10) {real, imag} */,
  {32'hc1d56f90, 32'h430cd4a8} /* (26, 28, 9) {real, imag} */,
  {32'h3f94b580, 32'hc180f63c} /* (26, 28, 8) {real, imag} */,
  {32'h431125f0, 32'h42005a54} /* (26, 28, 7) {real, imag} */,
  {32'h42b8c25b, 32'hc334c8e8} /* (26, 28, 6) {real, imag} */,
  {32'h423fdaf3, 32'h42851dee} /* (26, 28, 5) {real, imag} */,
  {32'h42699df1, 32'h41a6ceb6} /* (26, 28, 4) {real, imag} */,
  {32'h42a140f4, 32'h43352b96} /* (26, 28, 3) {real, imag} */,
  {32'hc2d9a4bf, 32'hc307b51e} /* (26, 28, 2) {real, imag} */,
  {32'hc425bc40, 32'hc40c1cdf} /* (26, 28, 1) {real, imag} */,
  {32'hc4eecf4c, 32'h00000000} /* (26, 28, 0) {real, imag} */,
  {32'hc43c529a, 32'h43e5c2f2} /* (26, 27, 31) {real, imag} */,
  {32'hc313a65a, 32'h42da5524} /* (26, 27, 30) {real, imag} */,
  {32'h42e2b984, 32'h412ad4a4} /* (26, 27, 29) {real, imag} */,
  {32'hc1c6f309, 32'hc15f8a80} /* (26, 27, 28) {real, imag} */,
  {32'h41f74c48, 32'h42b7b664} /* (26, 27, 27) {real, imag} */,
  {32'h431e479a, 32'h43177a5a} /* (26, 27, 26) {real, imag} */,
  {32'h421b15cb, 32'h3fad8b40} /* (26, 27, 25) {real, imag} */,
  {32'h4231cac1, 32'hc3323976} /* (26, 27, 24) {real, imag} */,
  {32'h40ae6fd4, 32'hc2d1a580} /* (26, 27, 23) {real, imag} */,
  {32'h414f34b0, 32'h423d8faf} /* (26, 27, 22) {real, imag} */,
  {32'hc2d86e72, 32'hc21c69d7} /* (26, 27, 21) {real, imag} */,
  {32'h42dafc12, 32'h418c0c58} /* (26, 27, 20) {real, imag} */,
  {32'hc259a958, 32'h42c2b90c} /* (26, 27, 19) {real, imag} */,
  {32'h41c735ee, 32'h4273bbaa} /* (26, 27, 18) {real, imag} */,
  {32'hc27b86b1, 32'hc2a40bb7} /* (26, 27, 17) {real, imag} */,
  {32'h42623b68, 32'h00000000} /* (26, 27, 16) {real, imag} */,
  {32'hc27b86b1, 32'h42a40bb7} /* (26, 27, 15) {real, imag} */,
  {32'h41c735ee, 32'hc273bbaa} /* (26, 27, 14) {real, imag} */,
  {32'hc259a958, 32'hc2c2b90c} /* (26, 27, 13) {real, imag} */,
  {32'h42dafc12, 32'hc18c0c58} /* (26, 27, 12) {real, imag} */,
  {32'hc2d86e72, 32'h421c69d7} /* (26, 27, 11) {real, imag} */,
  {32'h414f34b0, 32'hc23d8faf} /* (26, 27, 10) {real, imag} */,
  {32'h40ae6fd4, 32'h42d1a580} /* (26, 27, 9) {real, imag} */,
  {32'h4231cac1, 32'h43323976} /* (26, 27, 8) {real, imag} */,
  {32'h421b15cb, 32'hbfad8b40} /* (26, 27, 7) {real, imag} */,
  {32'h431e479a, 32'hc3177a5a} /* (26, 27, 6) {real, imag} */,
  {32'h41f74c48, 32'hc2b7b664} /* (26, 27, 5) {real, imag} */,
  {32'hc1c6f309, 32'h415f8a80} /* (26, 27, 4) {real, imag} */,
  {32'h42e2b984, 32'hc12ad4a4} /* (26, 27, 3) {real, imag} */,
  {32'hc313a65a, 32'hc2da5524} /* (26, 27, 2) {real, imag} */,
  {32'hc43c529a, 32'hc3e5c2f2} /* (26, 27, 1) {real, imag} */,
  {32'hc4e29bb5, 32'h00000000} /* (26, 27, 0) {real, imag} */,
  {32'hc4451256, 32'h43b50864} /* (26, 26, 31) {real, imag} */,
  {32'hc3087b43, 32'h43392f52} /* (26, 26, 30) {real, imag} */,
  {32'hc224ee06, 32'h427185ec} /* (26, 26, 29) {real, imag} */,
  {32'h42401906, 32'hc236ec02} /* (26, 26, 28) {real, imag} */,
  {32'hc164b126, 32'hc29f9d33} /* (26, 26, 27) {real, imag} */,
  {32'hc0a5323e, 32'hc1c05444} /* (26, 26, 26) {real, imag} */,
  {32'h419a4609, 32'hc274bf63} /* (26, 26, 25) {real, imag} */,
  {32'h40edbd92, 32'hc2577b8b} /* (26, 26, 24) {real, imag} */,
  {32'hc2d71b93, 32'h413838d8} /* (26, 26, 23) {real, imag} */,
  {32'h3f9ca450, 32'hc2732ffe} /* (26, 26, 22) {real, imag} */,
  {32'hc1d14bd2, 32'hc21f0bf0} /* (26, 26, 21) {real, imag} */,
  {32'h4214918e, 32'hc28dc008} /* (26, 26, 20) {real, imag} */,
  {32'h40e90af3, 32'h41a302cc} /* (26, 26, 19) {real, imag} */,
  {32'h4297cde1, 32'hc271ec02} /* (26, 26, 18) {real, imag} */,
  {32'h4248e643, 32'h4288c817} /* (26, 26, 17) {real, imag} */,
  {32'hc202dc58, 32'h00000000} /* (26, 26, 16) {real, imag} */,
  {32'h4248e643, 32'hc288c817} /* (26, 26, 15) {real, imag} */,
  {32'h4297cde1, 32'h4271ec02} /* (26, 26, 14) {real, imag} */,
  {32'h40e90af3, 32'hc1a302cc} /* (26, 26, 13) {real, imag} */,
  {32'h4214918e, 32'h428dc008} /* (26, 26, 12) {real, imag} */,
  {32'hc1d14bd2, 32'h421f0bf0} /* (26, 26, 11) {real, imag} */,
  {32'h3f9ca450, 32'h42732ffe} /* (26, 26, 10) {real, imag} */,
  {32'hc2d71b93, 32'hc13838d8} /* (26, 26, 9) {real, imag} */,
  {32'h40edbd92, 32'h42577b8b} /* (26, 26, 8) {real, imag} */,
  {32'h419a4609, 32'h4274bf63} /* (26, 26, 7) {real, imag} */,
  {32'hc0a5323e, 32'h41c05444} /* (26, 26, 6) {real, imag} */,
  {32'hc164b126, 32'h429f9d33} /* (26, 26, 5) {real, imag} */,
  {32'h42401906, 32'h4236ec02} /* (26, 26, 4) {real, imag} */,
  {32'hc224ee06, 32'hc27185ec} /* (26, 26, 3) {real, imag} */,
  {32'hc3087b43, 32'hc3392f52} /* (26, 26, 2) {real, imag} */,
  {32'hc4451256, 32'hc3b50864} /* (26, 26, 1) {real, imag} */,
  {32'hc4fbdf3c, 32'h00000000} /* (26, 26, 0) {real, imag} */,
  {32'hc4440b99, 32'h43a0a578} /* (26, 25, 31) {real, imag} */,
  {32'hc310635c, 32'h435cb938} /* (26, 25, 30) {real, imag} */,
  {32'hc0e770a0, 32'hc2632145} /* (26, 25, 29) {real, imag} */,
  {32'hc1d4619e, 32'hc28d68c9} /* (26, 25, 28) {real, imag} */,
  {32'h41e43796, 32'h423d682e} /* (26, 25, 27) {real, imag} */,
  {32'hc1fb93ad, 32'h4181a77e} /* (26, 25, 26) {real, imag} */,
  {32'h41f99534, 32'h402b26c0} /* (26, 25, 25) {real, imag} */,
  {32'h431c8590, 32'h421eb82a} /* (26, 25, 24) {real, imag} */,
  {32'hc21f0791, 32'h42047680} /* (26, 25, 23) {real, imag} */,
  {32'h42f1535f, 32'hc19a2939} /* (26, 25, 22) {real, imag} */,
  {32'hc24bd5a7, 32'hc1e9e9f0} /* (26, 25, 21) {real, imag} */,
  {32'h4194070d, 32'hc190c1a5} /* (26, 25, 20) {real, imag} */,
  {32'h41ad2dcf, 32'hc2488322} /* (26, 25, 19) {real, imag} */,
  {32'h4133e618, 32'h410d63d2} /* (26, 25, 18) {real, imag} */,
  {32'hc27722ca, 32'hc29f573c} /* (26, 25, 17) {real, imag} */,
  {32'h4086b3f0, 32'h00000000} /* (26, 25, 16) {real, imag} */,
  {32'hc27722ca, 32'h429f573c} /* (26, 25, 15) {real, imag} */,
  {32'h4133e618, 32'hc10d63d2} /* (26, 25, 14) {real, imag} */,
  {32'h41ad2dcf, 32'h42488322} /* (26, 25, 13) {real, imag} */,
  {32'h4194070d, 32'h4190c1a5} /* (26, 25, 12) {real, imag} */,
  {32'hc24bd5a7, 32'h41e9e9f0} /* (26, 25, 11) {real, imag} */,
  {32'h42f1535f, 32'h419a2939} /* (26, 25, 10) {real, imag} */,
  {32'hc21f0791, 32'hc2047680} /* (26, 25, 9) {real, imag} */,
  {32'h431c8590, 32'hc21eb82a} /* (26, 25, 8) {real, imag} */,
  {32'h41f99534, 32'hc02b26c0} /* (26, 25, 7) {real, imag} */,
  {32'hc1fb93ad, 32'hc181a77e} /* (26, 25, 6) {real, imag} */,
  {32'h41e43796, 32'hc23d682e} /* (26, 25, 5) {real, imag} */,
  {32'hc1d4619e, 32'h428d68c9} /* (26, 25, 4) {real, imag} */,
  {32'hc0e770a0, 32'h42632145} /* (26, 25, 3) {real, imag} */,
  {32'hc310635c, 32'hc35cb938} /* (26, 25, 2) {real, imag} */,
  {32'hc4440b99, 32'hc3a0a578} /* (26, 25, 1) {real, imag} */,
  {32'hc4c9bf53, 32'h00000000} /* (26, 25, 0) {real, imag} */,
  {32'hc437897a, 32'h430a6e54} /* (26, 24, 31) {real, imag} */,
  {32'hc2d806de, 32'h418ffe18} /* (26, 24, 30) {real, imag} */,
  {32'hc103ca00, 32'hc3115f28} /* (26, 24, 29) {real, imag} */,
  {32'h42da7bd0, 32'hbf982300} /* (26, 24, 28) {real, imag} */,
  {32'h41c5bdc8, 32'h432cb779} /* (26, 24, 27) {real, imag} */,
  {32'hc3240640, 32'hc26b47d3} /* (26, 24, 26) {real, imag} */,
  {32'h4252f18c, 32'h4258fe56} /* (26, 24, 25) {real, imag} */,
  {32'hc2802810, 32'h41692986} /* (26, 24, 24) {real, imag} */,
  {32'hc1c5fadd, 32'hc2c50628} /* (26, 24, 23) {real, imag} */,
  {32'hc0e8f010, 32'h41db0251} /* (26, 24, 22) {real, imag} */,
  {32'h40746390, 32'h4246273c} /* (26, 24, 21) {real, imag} */,
  {32'h42e76f38, 32'h4053b8b0} /* (26, 24, 20) {real, imag} */,
  {32'h419725eb, 32'hc203a6d7} /* (26, 24, 19) {real, imag} */,
  {32'hc24dd33c, 32'hc2e4c397} /* (26, 24, 18) {real, imag} */,
  {32'hc28d78de, 32'h42a9856b} /* (26, 24, 17) {real, imag} */,
  {32'hc228f64c, 32'h00000000} /* (26, 24, 16) {real, imag} */,
  {32'hc28d78de, 32'hc2a9856b} /* (26, 24, 15) {real, imag} */,
  {32'hc24dd33c, 32'h42e4c397} /* (26, 24, 14) {real, imag} */,
  {32'h419725eb, 32'h4203a6d7} /* (26, 24, 13) {real, imag} */,
  {32'h42e76f38, 32'hc053b8b0} /* (26, 24, 12) {real, imag} */,
  {32'h40746390, 32'hc246273c} /* (26, 24, 11) {real, imag} */,
  {32'hc0e8f010, 32'hc1db0251} /* (26, 24, 10) {real, imag} */,
  {32'hc1c5fadd, 32'h42c50628} /* (26, 24, 9) {real, imag} */,
  {32'hc2802810, 32'hc1692986} /* (26, 24, 8) {real, imag} */,
  {32'h4252f18c, 32'hc258fe56} /* (26, 24, 7) {real, imag} */,
  {32'hc3240640, 32'h426b47d3} /* (26, 24, 6) {real, imag} */,
  {32'h41c5bdc8, 32'hc32cb779} /* (26, 24, 5) {real, imag} */,
  {32'h42da7bd0, 32'h3f982300} /* (26, 24, 4) {real, imag} */,
  {32'hc103ca00, 32'h43115f28} /* (26, 24, 3) {real, imag} */,
  {32'hc2d806de, 32'hc18ffe18} /* (26, 24, 2) {real, imag} */,
  {32'hc437897a, 32'hc30a6e54} /* (26, 24, 1) {real, imag} */,
  {32'hc4a13e26, 32'h00000000} /* (26, 24, 0) {real, imag} */,
  {32'hc4380274, 32'h43053868} /* (26, 23, 31) {real, imag} */,
  {32'h41a14518, 32'hc1c15e34} /* (26, 23, 30) {real, imag} */,
  {32'h41552e80, 32'hc28e6558} /* (26, 23, 29) {real, imag} */,
  {32'h42dba475, 32'hc0f1cfb4} /* (26, 23, 28) {real, imag} */,
  {32'hc227cafd, 32'h4385bd65} /* (26, 23, 27) {real, imag} */,
  {32'hc222ca6e, 32'hc1a8ec36} /* (26, 23, 26) {real, imag} */,
  {32'hc1914228, 32'h41d5cc94} /* (26, 23, 25) {real, imag} */,
  {32'hc2cb48b4, 32'hc3071056} /* (26, 23, 24) {real, imag} */,
  {32'hc1a3e03c, 32'hbf5e49d8} /* (26, 23, 23) {real, imag} */,
  {32'hc23d3b58, 32'h423c4000} /* (26, 23, 22) {real, imag} */,
  {32'hc206478f, 32'h424813f2} /* (26, 23, 21) {real, imag} */,
  {32'h4040056c, 32'hc1ccdf9d} /* (26, 23, 20) {real, imag} */,
  {32'h42a72df1, 32'h3d5b1200} /* (26, 23, 19) {real, imag} */,
  {32'hc2bdffc7, 32'hc22283d0} /* (26, 23, 18) {real, imag} */,
  {32'h427f52f8, 32'hc09737f6} /* (26, 23, 17) {real, imag} */,
  {32'hc22ea0f0, 32'h00000000} /* (26, 23, 16) {real, imag} */,
  {32'h427f52f8, 32'h409737f6} /* (26, 23, 15) {real, imag} */,
  {32'hc2bdffc7, 32'h422283d0} /* (26, 23, 14) {real, imag} */,
  {32'h42a72df1, 32'hbd5b1200} /* (26, 23, 13) {real, imag} */,
  {32'h4040056c, 32'h41ccdf9d} /* (26, 23, 12) {real, imag} */,
  {32'hc206478f, 32'hc24813f2} /* (26, 23, 11) {real, imag} */,
  {32'hc23d3b58, 32'hc23c4000} /* (26, 23, 10) {real, imag} */,
  {32'hc1a3e03c, 32'h3f5e49d8} /* (26, 23, 9) {real, imag} */,
  {32'hc2cb48b4, 32'h43071056} /* (26, 23, 8) {real, imag} */,
  {32'hc1914228, 32'hc1d5cc94} /* (26, 23, 7) {real, imag} */,
  {32'hc222ca6e, 32'h41a8ec36} /* (26, 23, 6) {real, imag} */,
  {32'hc227cafd, 32'hc385bd65} /* (26, 23, 5) {real, imag} */,
  {32'h42dba475, 32'h40f1cfb4} /* (26, 23, 4) {real, imag} */,
  {32'h41552e80, 32'h428e6558} /* (26, 23, 3) {real, imag} */,
  {32'h41a14518, 32'h41c15e34} /* (26, 23, 2) {real, imag} */,
  {32'hc4380274, 32'hc3053868} /* (26, 23, 1) {real, imag} */,
  {32'hc48ad002, 32'h00000000} /* (26, 23, 0) {real, imag} */,
  {32'hc405fb36, 32'h438b8853} /* (26, 22, 31) {real, imag} */,
  {32'h4295af9d, 32'hc28832ca} /* (26, 22, 30) {real, imag} */,
  {32'h423655c2, 32'h4222eac4} /* (26, 22, 29) {real, imag} */,
  {32'h42e8303d, 32'hc19d1104} /* (26, 22, 28) {real, imag} */,
  {32'hc27a4ff6, 32'h4214eabe} /* (26, 22, 27) {real, imag} */,
  {32'h41523a70, 32'h42cf31b4} /* (26, 22, 26) {real, imag} */,
  {32'hc2a11ab8, 32'hc28c9bd4} /* (26, 22, 25) {real, imag} */,
  {32'hc299fbbd, 32'hc2559152} /* (26, 22, 24) {real, imag} */,
  {32'h42c5bdb5, 32'h42529b6c} /* (26, 22, 23) {real, imag} */,
  {32'hc135fc44, 32'hc22a21ca} /* (26, 22, 22) {real, imag} */,
  {32'h4119259c, 32'hc175c5d8} /* (26, 22, 21) {real, imag} */,
  {32'hc2553c76, 32'hc23e9c86} /* (26, 22, 20) {real, imag} */,
  {32'h419b3621, 32'h42921e73} /* (26, 22, 19) {real, imag} */,
  {32'hc14094ee, 32'h4208b1b8} /* (26, 22, 18) {real, imag} */,
  {32'hc1fb19cc, 32'hc22e139e} /* (26, 22, 17) {real, imag} */,
  {32'h422feff2, 32'h00000000} /* (26, 22, 16) {real, imag} */,
  {32'hc1fb19cc, 32'h422e139e} /* (26, 22, 15) {real, imag} */,
  {32'hc14094ee, 32'hc208b1b8} /* (26, 22, 14) {real, imag} */,
  {32'h419b3621, 32'hc2921e73} /* (26, 22, 13) {real, imag} */,
  {32'hc2553c76, 32'h423e9c86} /* (26, 22, 12) {real, imag} */,
  {32'h4119259c, 32'h4175c5d8} /* (26, 22, 11) {real, imag} */,
  {32'hc135fc44, 32'h422a21ca} /* (26, 22, 10) {real, imag} */,
  {32'h42c5bdb5, 32'hc2529b6c} /* (26, 22, 9) {real, imag} */,
  {32'hc299fbbd, 32'h42559152} /* (26, 22, 8) {real, imag} */,
  {32'hc2a11ab8, 32'h428c9bd4} /* (26, 22, 7) {real, imag} */,
  {32'h41523a70, 32'hc2cf31b4} /* (26, 22, 6) {real, imag} */,
  {32'hc27a4ff6, 32'hc214eabe} /* (26, 22, 5) {real, imag} */,
  {32'h42e8303d, 32'h419d1104} /* (26, 22, 4) {real, imag} */,
  {32'h423655c2, 32'hc222eac4} /* (26, 22, 3) {real, imag} */,
  {32'h4295af9d, 32'h428832ca} /* (26, 22, 2) {real, imag} */,
  {32'hc405fb36, 32'hc38b8853} /* (26, 22, 1) {real, imag} */,
  {32'hc3f01824, 32'h00000000} /* (26, 22, 0) {real, imag} */,
  {32'hc3cbdf6a, 32'h438fc76e} /* (26, 21, 31) {real, imag} */,
  {32'h4367fd9f, 32'h42ffa153} /* (26, 21, 30) {real, imag} */,
  {32'h41667e94, 32'h41b06dba} /* (26, 21, 29) {real, imag} */,
  {32'hc1cbe894, 32'hc295a00a} /* (26, 21, 28) {real, imag} */,
  {32'h425a5c5f, 32'hc24338be} /* (26, 21, 27) {real, imag} */,
  {32'h421ed5ef, 32'h4298050f} /* (26, 21, 26) {real, imag} */,
  {32'hc1bdbeba, 32'h40147b60} /* (26, 21, 25) {real, imag} */,
  {32'hc31d92a0, 32'h42b0ba1a} /* (26, 21, 24) {real, imag} */,
  {32'h400958b8, 32'hc2843f1e} /* (26, 21, 23) {real, imag} */,
  {32'h41f33632, 32'hc2957fce} /* (26, 21, 22) {real, imag} */,
  {32'h41407074, 32'h42e20958} /* (26, 21, 21) {real, imag} */,
  {32'h421b16ad, 32'hc22ce66a} /* (26, 21, 20) {real, imag} */,
  {32'hc19493e8, 32'hc0b91e44} /* (26, 21, 19) {real, imag} */,
  {32'h422c065e, 32'hc231e4cd} /* (26, 21, 18) {real, imag} */,
  {32'hc0bd3d0a, 32'h41b1f41e} /* (26, 21, 17) {real, imag} */,
  {32'h42d03896, 32'h00000000} /* (26, 21, 16) {real, imag} */,
  {32'hc0bd3d0a, 32'hc1b1f41e} /* (26, 21, 15) {real, imag} */,
  {32'h422c065e, 32'h4231e4cd} /* (26, 21, 14) {real, imag} */,
  {32'hc19493e8, 32'h40b91e44} /* (26, 21, 13) {real, imag} */,
  {32'h421b16ad, 32'h422ce66a} /* (26, 21, 12) {real, imag} */,
  {32'h41407074, 32'hc2e20958} /* (26, 21, 11) {real, imag} */,
  {32'h41f33632, 32'h42957fce} /* (26, 21, 10) {real, imag} */,
  {32'h400958b8, 32'h42843f1e} /* (26, 21, 9) {real, imag} */,
  {32'hc31d92a0, 32'hc2b0ba1a} /* (26, 21, 8) {real, imag} */,
  {32'hc1bdbeba, 32'hc0147b60} /* (26, 21, 7) {real, imag} */,
  {32'h421ed5ef, 32'hc298050f} /* (26, 21, 6) {real, imag} */,
  {32'h425a5c5f, 32'h424338be} /* (26, 21, 5) {real, imag} */,
  {32'hc1cbe894, 32'h4295a00a} /* (26, 21, 4) {real, imag} */,
  {32'h41667e94, 32'hc1b06dba} /* (26, 21, 3) {real, imag} */,
  {32'h4367fd9f, 32'hc2ffa153} /* (26, 21, 2) {real, imag} */,
  {32'hc3cbdf6a, 32'hc38fc76e} /* (26, 21, 1) {real, imag} */,
  {32'hc3a2f3fe, 32'h00000000} /* (26, 21, 0) {real, imag} */,
  {32'hc39fbed2, 32'hc105ede4} /* (26, 20, 31) {real, imag} */,
  {32'h4340896c, 32'hc1d908e9} /* (26, 20, 30) {real, imag} */,
  {32'h422e3511, 32'hc2992766} /* (26, 20, 29) {real, imag} */,
  {32'h428a5fac, 32'hc2bf372d} /* (26, 20, 28) {real, imag} */,
  {32'hc28042d3, 32'h429aa6ad} /* (26, 20, 27) {real, imag} */,
  {32'hc28719f6, 32'h42a1ce6e} /* (26, 20, 26) {real, imag} */,
  {32'h4063c1f0, 32'hc28bd2a8} /* (26, 20, 25) {real, imag} */,
  {32'h426516f9, 32'hc25c0780} /* (26, 20, 24) {real, imag} */,
  {32'h41970562, 32'h40e8e280} /* (26, 20, 23) {real, imag} */,
  {32'hc12c9ece, 32'hc0f4a1b8} /* (26, 20, 22) {real, imag} */,
  {32'h415d51ce, 32'hc1297863} /* (26, 20, 21) {real, imag} */,
  {32'hc1efcfbd, 32'hc117dd8c} /* (26, 20, 20) {real, imag} */,
  {32'hc2ccbf10, 32'h421f2119} /* (26, 20, 19) {real, imag} */,
  {32'h3e973ec0, 32'hc157d766} /* (26, 20, 18) {real, imag} */,
  {32'h41bdc3bc, 32'h411df496} /* (26, 20, 17) {real, imag} */,
  {32'h4268ca20, 32'h00000000} /* (26, 20, 16) {real, imag} */,
  {32'h41bdc3bc, 32'hc11df496} /* (26, 20, 15) {real, imag} */,
  {32'h3e973ec0, 32'h4157d766} /* (26, 20, 14) {real, imag} */,
  {32'hc2ccbf10, 32'hc21f2119} /* (26, 20, 13) {real, imag} */,
  {32'hc1efcfbd, 32'h4117dd8c} /* (26, 20, 12) {real, imag} */,
  {32'h415d51ce, 32'h41297863} /* (26, 20, 11) {real, imag} */,
  {32'hc12c9ece, 32'h40f4a1b8} /* (26, 20, 10) {real, imag} */,
  {32'h41970562, 32'hc0e8e280} /* (26, 20, 9) {real, imag} */,
  {32'h426516f9, 32'h425c0780} /* (26, 20, 8) {real, imag} */,
  {32'h4063c1f0, 32'h428bd2a8} /* (26, 20, 7) {real, imag} */,
  {32'hc28719f6, 32'hc2a1ce6e} /* (26, 20, 6) {real, imag} */,
  {32'hc28042d3, 32'hc29aa6ad} /* (26, 20, 5) {real, imag} */,
  {32'h428a5fac, 32'h42bf372d} /* (26, 20, 4) {real, imag} */,
  {32'h422e3511, 32'h42992766} /* (26, 20, 3) {real, imag} */,
  {32'h4340896c, 32'h41d908e9} /* (26, 20, 2) {real, imag} */,
  {32'hc39fbed2, 32'h4105ede4} /* (26, 20, 1) {real, imag} */,
  {32'hc38c6a42, 32'h00000000} /* (26, 20, 0) {real, imag} */,
  {32'hc37f8a12, 32'h421ebac2} /* (26, 19, 31) {real, imag} */,
  {32'h430a1430, 32'hc342db7a} /* (26, 19, 30) {real, imag} */,
  {32'h4269c5dc, 32'hc228fde8} /* (26, 19, 29) {real, imag} */,
  {32'h43292aed, 32'hc288701a} /* (26, 19, 28) {real, imag} */,
  {32'h41698a38, 32'h4286ff4e} /* (26, 19, 27) {real, imag} */,
  {32'h42448a58, 32'hc13d4914} /* (26, 19, 26) {real, imag} */,
  {32'hc2959086, 32'h424d5e46} /* (26, 19, 25) {real, imag} */,
  {32'h419845d2, 32'hc2c03baa} /* (26, 19, 24) {real, imag} */,
  {32'hc2c78ca6, 32'h423397b4} /* (26, 19, 23) {real, imag} */,
  {32'h41b7c73e, 32'hc251a0d8} /* (26, 19, 22) {real, imag} */,
  {32'hc2500e62, 32'hc1e3db68} /* (26, 19, 21) {real, imag} */,
  {32'h42783dce, 32'h40e8e016} /* (26, 19, 20) {real, imag} */,
  {32'hc2c6d3a2, 32'h42c24de8} /* (26, 19, 19) {real, imag} */,
  {32'h42295d1a, 32'h423e51f0} /* (26, 19, 18) {real, imag} */,
  {32'h40abcac0, 32'h4196274f} /* (26, 19, 17) {real, imag} */,
  {32'h420b7f9c, 32'h00000000} /* (26, 19, 16) {real, imag} */,
  {32'h40abcac0, 32'hc196274f} /* (26, 19, 15) {real, imag} */,
  {32'h42295d1a, 32'hc23e51f0} /* (26, 19, 14) {real, imag} */,
  {32'hc2c6d3a2, 32'hc2c24de8} /* (26, 19, 13) {real, imag} */,
  {32'h42783dce, 32'hc0e8e016} /* (26, 19, 12) {real, imag} */,
  {32'hc2500e62, 32'h41e3db68} /* (26, 19, 11) {real, imag} */,
  {32'h41b7c73e, 32'h4251a0d8} /* (26, 19, 10) {real, imag} */,
  {32'hc2c78ca6, 32'hc23397b4} /* (26, 19, 9) {real, imag} */,
  {32'h419845d2, 32'h42c03baa} /* (26, 19, 8) {real, imag} */,
  {32'hc2959086, 32'hc24d5e46} /* (26, 19, 7) {real, imag} */,
  {32'h42448a58, 32'h413d4914} /* (26, 19, 6) {real, imag} */,
  {32'h41698a38, 32'hc286ff4e} /* (26, 19, 5) {real, imag} */,
  {32'h43292aed, 32'h4288701a} /* (26, 19, 4) {real, imag} */,
  {32'h4269c5dc, 32'h4228fde8} /* (26, 19, 3) {real, imag} */,
  {32'h430a1430, 32'h4342db7a} /* (26, 19, 2) {real, imag} */,
  {32'hc37f8a12, 32'hc21ebac2} /* (26, 19, 1) {real, imag} */,
  {32'hc24f2cce, 32'h00000000} /* (26, 19, 0) {real, imag} */,
  {32'hc14b41b0, 32'h4315b7b6} /* (26, 18, 31) {real, imag} */,
  {32'h432f5602, 32'hc325420a} /* (26, 18, 30) {real, imag} */,
  {32'h4061a0f8, 32'hc302bf5c} /* (26, 18, 29) {real, imag} */,
  {32'h42ee0968, 32'h41d1b17e} /* (26, 18, 28) {real, imag} */,
  {32'h41a3406a, 32'h41888484} /* (26, 18, 27) {real, imag} */,
  {32'h42e96b2d, 32'hc2afb8c4} /* (26, 18, 26) {real, imag} */,
  {32'hc2b15c77, 32'h42d5b624} /* (26, 18, 25) {real, imag} */,
  {32'hc27a6935, 32'hc1108ba8} /* (26, 18, 24) {real, imag} */,
  {32'h41e6c070, 32'h416a5ea5} /* (26, 18, 23) {real, imag} */,
  {32'hc28abc54, 32'hc0da53a0} /* (26, 18, 22) {real, imag} */,
  {32'hc288c2c6, 32'hc2aea71e} /* (26, 18, 21) {real, imag} */,
  {32'hc11016c2, 32'hc16744ca} /* (26, 18, 20) {real, imag} */,
  {32'hc20cf760, 32'hc23a52a4} /* (26, 18, 19) {real, imag} */,
  {32'hc272cfc0, 32'h41928647} /* (26, 18, 18) {real, imag} */,
  {32'h41792552, 32'h4045c9d8} /* (26, 18, 17) {real, imag} */,
  {32'hc23dba8c, 32'h00000000} /* (26, 18, 16) {real, imag} */,
  {32'h41792552, 32'hc045c9d8} /* (26, 18, 15) {real, imag} */,
  {32'hc272cfc0, 32'hc1928647} /* (26, 18, 14) {real, imag} */,
  {32'hc20cf760, 32'h423a52a4} /* (26, 18, 13) {real, imag} */,
  {32'hc11016c2, 32'h416744ca} /* (26, 18, 12) {real, imag} */,
  {32'hc288c2c6, 32'h42aea71e} /* (26, 18, 11) {real, imag} */,
  {32'hc28abc54, 32'h40da53a0} /* (26, 18, 10) {real, imag} */,
  {32'h41e6c070, 32'hc16a5ea5} /* (26, 18, 9) {real, imag} */,
  {32'hc27a6935, 32'h41108ba8} /* (26, 18, 8) {real, imag} */,
  {32'hc2b15c77, 32'hc2d5b624} /* (26, 18, 7) {real, imag} */,
  {32'h42e96b2d, 32'h42afb8c4} /* (26, 18, 6) {real, imag} */,
  {32'h41a3406a, 32'hc1888484} /* (26, 18, 5) {real, imag} */,
  {32'h42ee0968, 32'hc1d1b17e} /* (26, 18, 4) {real, imag} */,
  {32'h4061a0f8, 32'h4302bf5c} /* (26, 18, 3) {real, imag} */,
  {32'h432f5602, 32'h4325420a} /* (26, 18, 2) {real, imag} */,
  {32'hc14b41b0, 32'hc315b7b6} /* (26, 18, 1) {real, imag} */,
  {32'h42124940, 32'h00000000} /* (26, 18, 0) {real, imag} */,
  {32'h42647b58, 32'h4343adac} /* (26, 17, 31) {real, imag} */,
  {32'h4248a97f, 32'hc2ca7066} /* (26, 17, 30) {real, imag} */,
  {32'hc31130d5, 32'hc3130cce} /* (26, 17, 29) {real, imag} */,
  {32'h43152bb8, 32'h40960ac4} /* (26, 17, 28) {real, imag} */,
  {32'h41a0caf9, 32'hc0b6a2cc} /* (26, 17, 27) {real, imag} */,
  {32'h42953445, 32'hc170c04c} /* (26, 17, 26) {real, imag} */,
  {32'h408a16d0, 32'hc0e89448} /* (26, 17, 25) {real, imag} */,
  {32'hc2b4ecd0, 32'hc1e9721c} /* (26, 17, 24) {real, imag} */,
  {32'h42945ab2, 32'h4203d34d} /* (26, 17, 23) {real, imag} */,
  {32'h427288b1, 32'h426591ea} /* (26, 17, 22) {real, imag} */,
  {32'h4298cb4e, 32'h413a5f56} /* (26, 17, 21) {real, imag} */,
  {32'hc2555128, 32'h41893337} /* (26, 17, 20) {real, imag} */,
  {32'hc29d735a, 32'hc2cb502b} /* (26, 17, 19) {real, imag} */,
  {32'hc2869f82, 32'hc0cebf80} /* (26, 17, 18) {real, imag} */,
  {32'hc1db0d09, 32'h41d38be8} /* (26, 17, 17) {real, imag} */,
  {32'h41ab6994, 32'h00000000} /* (26, 17, 16) {real, imag} */,
  {32'hc1db0d09, 32'hc1d38be8} /* (26, 17, 15) {real, imag} */,
  {32'hc2869f82, 32'h40cebf80} /* (26, 17, 14) {real, imag} */,
  {32'hc29d735a, 32'h42cb502b} /* (26, 17, 13) {real, imag} */,
  {32'hc2555128, 32'hc1893337} /* (26, 17, 12) {real, imag} */,
  {32'h4298cb4e, 32'hc13a5f56} /* (26, 17, 11) {real, imag} */,
  {32'h427288b1, 32'hc26591ea} /* (26, 17, 10) {real, imag} */,
  {32'h42945ab2, 32'hc203d34d} /* (26, 17, 9) {real, imag} */,
  {32'hc2b4ecd0, 32'h41e9721c} /* (26, 17, 8) {real, imag} */,
  {32'h408a16d0, 32'h40e89448} /* (26, 17, 7) {real, imag} */,
  {32'h42953445, 32'h4170c04c} /* (26, 17, 6) {real, imag} */,
  {32'h41a0caf9, 32'h40b6a2cc} /* (26, 17, 5) {real, imag} */,
  {32'h43152bb8, 32'hc0960ac4} /* (26, 17, 4) {real, imag} */,
  {32'hc31130d5, 32'h43130cce} /* (26, 17, 3) {real, imag} */,
  {32'h4248a97f, 32'h42ca7066} /* (26, 17, 2) {real, imag} */,
  {32'h42647b58, 32'hc343adac} /* (26, 17, 1) {real, imag} */,
  {32'h42a99c52, 32'h00000000} /* (26, 17, 0) {real, imag} */,
  {32'h431d8860, 32'h434c6e82} /* (26, 16, 31) {real, imag} */,
  {32'hc0ad04b0, 32'hc2756e20} /* (26, 16, 30) {real, imag} */,
  {32'hc22cf7f8, 32'hc300fcbc} /* (26, 16, 29) {real, imag} */,
  {32'h41c5a3b4, 32'hc20f5bba} /* (26, 16, 28) {real, imag} */,
  {32'h423570c9, 32'hc28aee3a} /* (26, 16, 27) {real, imag} */,
  {32'h410db194, 32'h428047bb} /* (26, 16, 26) {real, imag} */,
  {32'h4197ab59, 32'h42c15680} /* (26, 16, 25) {real, imag} */,
  {32'h41d0ae6e, 32'hc112b786} /* (26, 16, 24) {real, imag} */,
  {32'h4141b806, 32'h40836bb0} /* (26, 16, 23) {real, imag} */,
  {32'h42988820, 32'hc1b2472a} /* (26, 16, 22) {real, imag} */,
  {32'h42b289e6, 32'h42d5ab21} /* (26, 16, 21) {real, imag} */,
  {32'hc271a44a, 32'hc222561c} /* (26, 16, 20) {real, imag} */,
  {32'h4019faf8, 32'hc1107d02} /* (26, 16, 19) {real, imag} */,
  {32'h424e9afd, 32'h42b64ef2} /* (26, 16, 18) {real, imag} */,
  {32'hc19b73da, 32'hc1c0b847} /* (26, 16, 17) {real, imag} */,
  {32'h42bc5798, 32'h00000000} /* (26, 16, 16) {real, imag} */,
  {32'hc19b73da, 32'h41c0b847} /* (26, 16, 15) {real, imag} */,
  {32'h424e9afd, 32'hc2b64ef2} /* (26, 16, 14) {real, imag} */,
  {32'h4019faf8, 32'h41107d02} /* (26, 16, 13) {real, imag} */,
  {32'hc271a44a, 32'h4222561c} /* (26, 16, 12) {real, imag} */,
  {32'h42b289e6, 32'hc2d5ab21} /* (26, 16, 11) {real, imag} */,
  {32'h42988820, 32'h41b2472a} /* (26, 16, 10) {real, imag} */,
  {32'h4141b806, 32'hc0836bb0} /* (26, 16, 9) {real, imag} */,
  {32'h41d0ae6e, 32'h4112b786} /* (26, 16, 8) {real, imag} */,
  {32'h4197ab59, 32'hc2c15680} /* (26, 16, 7) {real, imag} */,
  {32'h410db194, 32'hc28047bb} /* (26, 16, 6) {real, imag} */,
  {32'h423570c9, 32'h428aee3a} /* (26, 16, 5) {real, imag} */,
  {32'h41c5a3b4, 32'h420f5bba} /* (26, 16, 4) {real, imag} */,
  {32'hc22cf7f8, 32'h4300fcbc} /* (26, 16, 3) {real, imag} */,
  {32'hc0ad04b0, 32'h42756e20} /* (26, 16, 2) {real, imag} */,
  {32'h431d8860, 32'hc34c6e82} /* (26, 16, 1) {real, imag} */,
  {32'h432db864, 32'h00000000} /* (26, 16, 0) {real, imag} */,
  {32'h4353c446, 32'h430cc49c} /* (26, 15, 31) {real, imag} */,
  {32'hc24c3d65, 32'hc2c73f7e} /* (26, 15, 30) {real, imag} */,
  {32'h41365950, 32'h42b9d4d7} /* (26, 15, 29) {real, imag} */,
  {32'h410fa278, 32'hc244bf12} /* (26, 15, 28) {real, imag} */,
  {32'h428c0e8a, 32'hc0eac1a4} /* (26, 15, 27) {real, imag} */,
  {32'h42a92063, 32'h4229ca95} /* (26, 15, 26) {real, imag} */,
  {32'h4270e0d2, 32'h43013370} /* (26, 15, 25) {real, imag} */,
  {32'h43241da9, 32'hc2a0871b} /* (26, 15, 24) {real, imag} */,
  {32'hc2bba6b4, 32'hc28721fc} /* (26, 15, 23) {real, imag} */,
  {32'hc205615f, 32'hc1ec79f4} /* (26, 15, 22) {real, imag} */,
  {32'h41a4772e, 32'h428644a9} /* (26, 15, 21) {real, imag} */,
  {32'hc1889228, 32'hc24d0a1a} /* (26, 15, 20) {real, imag} */,
  {32'hc3301e23, 32'h42589dc2} /* (26, 15, 19) {real, imag} */,
  {32'h41581fc0, 32'h42297097} /* (26, 15, 18) {real, imag} */,
  {32'h41b296cb, 32'h4220d368} /* (26, 15, 17) {real, imag} */,
  {32'h42b44be2, 32'h00000000} /* (26, 15, 16) {real, imag} */,
  {32'h41b296cb, 32'hc220d368} /* (26, 15, 15) {real, imag} */,
  {32'h41581fc0, 32'hc2297097} /* (26, 15, 14) {real, imag} */,
  {32'hc3301e23, 32'hc2589dc2} /* (26, 15, 13) {real, imag} */,
  {32'hc1889228, 32'h424d0a1a} /* (26, 15, 12) {real, imag} */,
  {32'h41a4772e, 32'hc28644a9} /* (26, 15, 11) {real, imag} */,
  {32'hc205615f, 32'h41ec79f4} /* (26, 15, 10) {real, imag} */,
  {32'hc2bba6b4, 32'h428721fc} /* (26, 15, 9) {real, imag} */,
  {32'h43241da9, 32'h42a0871b} /* (26, 15, 8) {real, imag} */,
  {32'h4270e0d2, 32'hc3013370} /* (26, 15, 7) {real, imag} */,
  {32'h42a92063, 32'hc229ca95} /* (26, 15, 6) {real, imag} */,
  {32'h428c0e8a, 32'h40eac1a4} /* (26, 15, 5) {real, imag} */,
  {32'h410fa278, 32'h4244bf12} /* (26, 15, 4) {real, imag} */,
  {32'h41365950, 32'hc2b9d4d7} /* (26, 15, 3) {real, imag} */,
  {32'hc24c3d65, 32'h42c73f7e} /* (26, 15, 2) {real, imag} */,
  {32'h4353c446, 32'hc30cc49c} /* (26, 15, 1) {real, imag} */,
  {32'hc3937288, 32'h00000000} /* (26, 15, 0) {real, imag} */,
  {32'h433e7d7b, 32'h43673954} /* (26, 14, 31) {real, imag} */,
  {32'h4268618e, 32'h42929219} /* (26, 14, 30) {real, imag} */,
  {32'hc1c60bad, 32'h407b0fa0} /* (26, 14, 29) {real, imag} */,
  {32'hc1ca1f8a, 32'h41c97e1a} /* (26, 14, 28) {real, imag} */,
  {32'h425b351b, 32'hc101c81c} /* (26, 14, 27) {real, imag} */,
  {32'hc08988d0, 32'hc1b77048} /* (26, 14, 26) {real, imag} */,
  {32'h420e8450, 32'h3fef9100} /* (26, 14, 25) {real, imag} */,
  {32'h42a669c6, 32'hc30271f0} /* (26, 14, 24) {real, imag} */,
  {32'h4212424c, 32'hc10afd2d} /* (26, 14, 23) {real, imag} */,
  {32'h41d0d074, 32'h427e9b82} /* (26, 14, 22) {real, imag} */,
  {32'h4232c91d, 32'h4228a945} /* (26, 14, 21) {real, imag} */,
  {32'h4081a59c, 32'h40f094d4} /* (26, 14, 20) {real, imag} */,
  {32'hc29587fc, 32'hc13ef39a} /* (26, 14, 19) {real, imag} */,
  {32'hc293b698, 32'h42450170} /* (26, 14, 18) {real, imag} */,
  {32'hc0a05a71, 32'h42204b1a} /* (26, 14, 17) {real, imag} */,
  {32'h417dc03f, 32'h00000000} /* (26, 14, 16) {real, imag} */,
  {32'hc0a05a71, 32'hc2204b1a} /* (26, 14, 15) {real, imag} */,
  {32'hc293b698, 32'hc2450170} /* (26, 14, 14) {real, imag} */,
  {32'hc29587fc, 32'h413ef39a} /* (26, 14, 13) {real, imag} */,
  {32'h4081a59c, 32'hc0f094d4} /* (26, 14, 12) {real, imag} */,
  {32'h4232c91d, 32'hc228a945} /* (26, 14, 11) {real, imag} */,
  {32'h41d0d074, 32'hc27e9b82} /* (26, 14, 10) {real, imag} */,
  {32'h4212424c, 32'h410afd2d} /* (26, 14, 9) {real, imag} */,
  {32'h42a669c6, 32'h430271f0} /* (26, 14, 8) {real, imag} */,
  {32'h420e8450, 32'hbfef9100} /* (26, 14, 7) {real, imag} */,
  {32'hc08988d0, 32'h41b77048} /* (26, 14, 6) {real, imag} */,
  {32'h425b351b, 32'h4101c81c} /* (26, 14, 5) {real, imag} */,
  {32'hc1ca1f8a, 32'hc1c97e1a} /* (26, 14, 4) {real, imag} */,
  {32'hc1c60bad, 32'hc07b0fa0} /* (26, 14, 3) {real, imag} */,
  {32'h4268618e, 32'hc2929219} /* (26, 14, 2) {real, imag} */,
  {32'h433e7d7b, 32'hc3673954} /* (26, 14, 1) {real, imag} */,
  {32'hc3a19fc0, 32'h00000000} /* (26, 14, 0) {real, imag} */,
  {32'h435df242, 32'h43423cd0} /* (26, 13, 31) {real, imag} */,
  {32'hc220cd76, 32'h4200f428} /* (26, 13, 30) {real, imag} */,
  {32'hc16bb8b2, 32'hc2850a23} /* (26, 13, 29) {real, imag} */,
  {32'hc2e948de, 32'h430f5740} /* (26, 13, 28) {real, imag} */,
  {32'h41c0d37e, 32'hc2cd44fa} /* (26, 13, 27) {real, imag} */,
  {32'h421c167c, 32'hc1ff7172} /* (26, 13, 26) {real, imag} */,
  {32'h430d7a31, 32'hc295c476} /* (26, 13, 25) {real, imag} */,
  {32'h423383b5, 32'hc25c180c} /* (26, 13, 24) {real, imag} */,
  {32'hc220b768, 32'hc0ab0d7c} /* (26, 13, 23) {real, imag} */,
  {32'hc1d90aea, 32'h41759550} /* (26, 13, 22) {real, imag} */,
  {32'h424e3c2a, 32'h4123e2df} /* (26, 13, 21) {real, imag} */,
  {32'hc1bb6e3c, 32'hc00aed24} /* (26, 13, 20) {real, imag} */,
  {32'h41a1703e, 32'h42819a84} /* (26, 13, 19) {real, imag} */,
  {32'h421ac416, 32'hc26bea44} /* (26, 13, 18) {real, imag} */,
  {32'hc2185eb2, 32'hc1d1228b} /* (26, 13, 17) {real, imag} */,
  {32'hc16fcb26, 32'h00000000} /* (26, 13, 16) {real, imag} */,
  {32'hc2185eb2, 32'h41d1228b} /* (26, 13, 15) {real, imag} */,
  {32'h421ac416, 32'h426bea44} /* (26, 13, 14) {real, imag} */,
  {32'h41a1703e, 32'hc2819a84} /* (26, 13, 13) {real, imag} */,
  {32'hc1bb6e3c, 32'h400aed24} /* (26, 13, 12) {real, imag} */,
  {32'h424e3c2a, 32'hc123e2df} /* (26, 13, 11) {real, imag} */,
  {32'hc1d90aea, 32'hc1759550} /* (26, 13, 10) {real, imag} */,
  {32'hc220b768, 32'h40ab0d7c} /* (26, 13, 9) {real, imag} */,
  {32'h423383b5, 32'h425c180c} /* (26, 13, 8) {real, imag} */,
  {32'h430d7a31, 32'h4295c476} /* (26, 13, 7) {real, imag} */,
  {32'h421c167c, 32'h41ff7172} /* (26, 13, 6) {real, imag} */,
  {32'h41c0d37e, 32'h42cd44fa} /* (26, 13, 5) {real, imag} */,
  {32'hc2e948de, 32'hc30f5740} /* (26, 13, 4) {real, imag} */,
  {32'hc16bb8b2, 32'h42850a23} /* (26, 13, 3) {real, imag} */,
  {32'hc220cd76, 32'hc200f428} /* (26, 13, 2) {real, imag} */,
  {32'h435df242, 32'hc3423cd0} /* (26, 13, 1) {real, imag} */,
  {32'hc3841026, 32'h00000000} /* (26, 13, 0) {real, imag} */,
  {32'h42bb3e40, 32'h428ac1dc} /* (26, 12, 31) {real, imag} */,
  {32'hc276f2ee, 32'hc288646e} /* (26, 12, 30) {real, imag} */,
  {32'h41ab3bc2, 32'hc272378c} /* (26, 12, 29) {real, imag} */,
  {32'hc1907da0, 32'hc2362d4e} /* (26, 12, 28) {real, imag} */,
  {32'hc23cb4e8, 32'hc2907989} /* (26, 12, 27) {real, imag} */,
  {32'h42801018, 32'h40ba9e78} /* (26, 12, 26) {real, imag} */,
  {32'h429c174c, 32'hc15bc4d0} /* (26, 12, 25) {real, imag} */,
  {32'hc1650664, 32'hbfc397f0} /* (26, 12, 24) {real, imag} */,
  {32'h41c7ba08, 32'hc21a1114} /* (26, 12, 23) {real, imag} */,
  {32'h41ec9caf, 32'h4072c930} /* (26, 12, 22) {real, imag} */,
  {32'h4258b178, 32'h40f6b3f2} /* (26, 12, 21) {real, imag} */,
  {32'h412b7a62, 32'hc27c283b} /* (26, 12, 20) {real, imag} */,
  {32'hc173fa38, 32'hc1ab5eea} /* (26, 12, 19) {real, imag} */,
  {32'h4249e820, 32'hc2191a68} /* (26, 12, 18) {real, imag} */,
  {32'h42c9f08d, 32'h422aa97e} /* (26, 12, 17) {real, imag} */,
  {32'h424a5922, 32'h00000000} /* (26, 12, 16) {real, imag} */,
  {32'h42c9f08d, 32'hc22aa97e} /* (26, 12, 15) {real, imag} */,
  {32'h4249e820, 32'h42191a68} /* (26, 12, 14) {real, imag} */,
  {32'hc173fa38, 32'h41ab5eea} /* (26, 12, 13) {real, imag} */,
  {32'h412b7a62, 32'h427c283b} /* (26, 12, 12) {real, imag} */,
  {32'h4258b178, 32'hc0f6b3f2} /* (26, 12, 11) {real, imag} */,
  {32'h41ec9caf, 32'hc072c930} /* (26, 12, 10) {real, imag} */,
  {32'h41c7ba08, 32'h421a1114} /* (26, 12, 9) {real, imag} */,
  {32'hc1650664, 32'h3fc397f0} /* (26, 12, 8) {real, imag} */,
  {32'h429c174c, 32'h415bc4d0} /* (26, 12, 7) {real, imag} */,
  {32'h42801018, 32'hc0ba9e78} /* (26, 12, 6) {real, imag} */,
  {32'hc23cb4e8, 32'h42907989} /* (26, 12, 5) {real, imag} */,
  {32'hc1907da0, 32'h42362d4e} /* (26, 12, 4) {real, imag} */,
  {32'h41ab3bc2, 32'h4272378c} /* (26, 12, 3) {real, imag} */,
  {32'hc276f2ee, 32'h4288646e} /* (26, 12, 2) {real, imag} */,
  {32'h42bb3e40, 32'hc28ac1dc} /* (26, 12, 1) {real, imag} */,
  {32'hc36eb1cc, 32'h00000000} /* (26, 12, 0) {real, imag} */,
  {32'hc1c46b68, 32'h431649e6} /* (26, 11, 31) {real, imag} */,
  {32'hc32f3e3d, 32'h428871c9} /* (26, 11, 30) {real, imag} */,
  {32'h4280b844, 32'hc301211d} /* (26, 11, 29) {real, imag} */,
  {32'h4312fbd2, 32'hc30139eb} /* (26, 11, 28) {real, imag} */,
  {32'hc2989d60, 32'hc1ce86a9} /* (26, 11, 27) {real, imag} */,
  {32'h424ede01, 32'hc202740e} /* (26, 11, 26) {real, imag} */,
  {32'hc228a45b, 32'hc29c3249} /* (26, 11, 25) {real, imag} */,
  {32'h4233cd4a, 32'hc1e5e19e} /* (26, 11, 24) {real, imag} */,
  {32'h414623f6, 32'hc1c94223} /* (26, 11, 23) {real, imag} */,
  {32'hc2def404, 32'h4280b214} /* (26, 11, 22) {real, imag} */,
  {32'hc1b34f22, 32'h4295244c} /* (26, 11, 21) {real, imag} */,
  {32'hc2a2495a, 32'hc12ff948} /* (26, 11, 20) {real, imag} */,
  {32'h428435de, 32'hc25d9cc4} /* (26, 11, 19) {real, imag} */,
  {32'hc1d06c5c, 32'hc2386107} /* (26, 11, 18) {real, imag} */,
  {32'h4133e401, 32'hc1a95bd6} /* (26, 11, 17) {real, imag} */,
  {32'h42054d00, 32'h00000000} /* (26, 11, 16) {real, imag} */,
  {32'h4133e401, 32'h41a95bd6} /* (26, 11, 15) {real, imag} */,
  {32'hc1d06c5c, 32'h42386107} /* (26, 11, 14) {real, imag} */,
  {32'h428435de, 32'h425d9cc4} /* (26, 11, 13) {real, imag} */,
  {32'hc2a2495a, 32'h412ff948} /* (26, 11, 12) {real, imag} */,
  {32'hc1b34f22, 32'hc295244c} /* (26, 11, 11) {real, imag} */,
  {32'hc2def404, 32'hc280b214} /* (26, 11, 10) {real, imag} */,
  {32'h414623f6, 32'h41c94223} /* (26, 11, 9) {real, imag} */,
  {32'h4233cd4a, 32'h41e5e19e} /* (26, 11, 8) {real, imag} */,
  {32'hc228a45b, 32'h429c3249} /* (26, 11, 7) {real, imag} */,
  {32'h424ede01, 32'h4202740e} /* (26, 11, 6) {real, imag} */,
  {32'hc2989d60, 32'h41ce86a9} /* (26, 11, 5) {real, imag} */,
  {32'h4312fbd2, 32'h430139eb} /* (26, 11, 4) {real, imag} */,
  {32'h4280b844, 32'h4301211d} /* (26, 11, 3) {real, imag} */,
  {32'hc32f3e3d, 32'hc28871c9} /* (26, 11, 2) {real, imag} */,
  {32'hc1c46b68, 32'hc31649e6} /* (26, 11, 1) {real, imag} */,
  {32'hc24ec1cc, 32'h00000000} /* (26, 11, 0) {real, imag} */,
  {32'h42bdbf90, 32'h438c0e45} /* (26, 10, 31) {real, imag} */,
  {32'hc31fbbda, 32'h42c5ee18} /* (26, 10, 30) {real, imag} */,
  {32'h41b66cfc, 32'hc287ac5e} /* (26, 10, 29) {real, imag} */,
  {32'h431c7470, 32'hc2d3b99b} /* (26, 10, 28) {real, imag} */,
  {32'h42524044, 32'h4123647e} /* (26, 10, 27) {real, imag} */,
  {32'h42976c56, 32'hc2151b94} /* (26, 10, 26) {real, imag} */,
  {32'h400f5480, 32'h423af489} /* (26, 10, 25) {real, imag} */,
  {32'h42cdfc1b, 32'hc204e488} /* (26, 10, 24) {real, imag} */,
  {32'hc311752a, 32'h4242a608} /* (26, 10, 23) {real, imag} */,
  {32'h429cf8c2, 32'h42d826d3} /* (26, 10, 22) {real, imag} */,
  {32'hc19d05e4, 32'h42d7832b} /* (26, 10, 21) {real, imag} */,
  {32'hc23275f2, 32'h42033994} /* (26, 10, 20) {real, imag} */,
  {32'h41b04d7b, 32'h42cc358f} /* (26, 10, 19) {real, imag} */,
  {32'h4251c4ac, 32'hc2791c1c} /* (26, 10, 18) {real, imag} */,
  {32'h405616c0, 32'h41c49fd4} /* (26, 10, 17) {real, imag} */,
  {32'h429e4a2b, 32'h00000000} /* (26, 10, 16) {real, imag} */,
  {32'h405616c0, 32'hc1c49fd4} /* (26, 10, 15) {real, imag} */,
  {32'h4251c4ac, 32'h42791c1c} /* (26, 10, 14) {real, imag} */,
  {32'h41b04d7b, 32'hc2cc358f} /* (26, 10, 13) {real, imag} */,
  {32'hc23275f2, 32'hc2033994} /* (26, 10, 12) {real, imag} */,
  {32'hc19d05e4, 32'hc2d7832b} /* (26, 10, 11) {real, imag} */,
  {32'h429cf8c2, 32'hc2d826d3} /* (26, 10, 10) {real, imag} */,
  {32'hc311752a, 32'hc242a608} /* (26, 10, 9) {real, imag} */,
  {32'h42cdfc1b, 32'h4204e488} /* (26, 10, 8) {real, imag} */,
  {32'h400f5480, 32'hc23af489} /* (26, 10, 7) {real, imag} */,
  {32'h42976c56, 32'h42151b94} /* (26, 10, 6) {real, imag} */,
  {32'h42524044, 32'hc123647e} /* (26, 10, 5) {real, imag} */,
  {32'h431c7470, 32'h42d3b99b} /* (26, 10, 4) {real, imag} */,
  {32'h41b66cfc, 32'h4287ac5e} /* (26, 10, 3) {real, imag} */,
  {32'hc31fbbda, 32'hc2c5ee18} /* (26, 10, 2) {real, imag} */,
  {32'h42bdbf90, 32'hc38c0e45} /* (26, 10, 1) {real, imag} */,
  {32'hc3670cb1, 32'h00000000} /* (26, 10, 0) {real, imag} */,
  {32'h4200fae0, 32'h43aaa79f} /* (26, 9, 31) {real, imag} */,
  {32'hc349e8c3, 32'h42e3576b} /* (26, 9, 30) {real, imag} */,
  {32'h423f8efe, 32'hc2bc90ac} /* (26, 9, 29) {real, imag} */,
  {32'h42c252f7, 32'hc28ba487} /* (26, 9, 28) {real, imag} */,
  {32'hc011dd30, 32'hbc2a8000} /* (26, 9, 27) {real, imag} */,
  {32'h3f9e7b30, 32'hc2562399} /* (26, 9, 26) {real, imag} */,
  {32'hc2af6dce, 32'h423f39a8} /* (26, 9, 25) {real, imag} */,
  {32'h407c5d10, 32'h418fd734} /* (26, 9, 24) {real, imag} */,
  {32'hc0ce7b4e, 32'hc1297a02} /* (26, 9, 23) {real, imag} */,
  {32'hc271d9ec, 32'h429c8ee4} /* (26, 9, 22) {real, imag} */,
  {32'h417dda74, 32'h410bafee} /* (26, 9, 21) {real, imag} */,
  {32'h41a3291c, 32'h41e47381} /* (26, 9, 20) {real, imag} */,
  {32'hc2c5f8df, 32'hc2566494} /* (26, 9, 19) {real, imag} */,
  {32'hc27c634a, 32'h40b43064} /* (26, 9, 18) {real, imag} */,
  {32'h40201c38, 32'h419480fc} /* (26, 9, 17) {real, imag} */,
  {32'h42c00884, 32'h00000000} /* (26, 9, 16) {real, imag} */,
  {32'h40201c38, 32'hc19480fc} /* (26, 9, 15) {real, imag} */,
  {32'hc27c634a, 32'hc0b43064} /* (26, 9, 14) {real, imag} */,
  {32'hc2c5f8df, 32'h42566494} /* (26, 9, 13) {real, imag} */,
  {32'h41a3291c, 32'hc1e47381} /* (26, 9, 12) {real, imag} */,
  {32'h417dda74, 32'hc10bafee} /* (26, 9, 11) {real, imag} */,
  {32'hc271d9ec, 32'hc29c8ee4} /* (26, 9, 10) {real, imag} */,
  {32'hc0ce7b4e, 32'h41297a02} /* (26, 9, 9) {real, imag} */,
  {32'h407c5d10, 32'hc18fd734} /* (26, 9, 8) {real, imag} */,
  {32'hc2af6dce, 32'hc23f39a8} /* (26, 9, 7) {real, imag} */,
  {32'h3f9e7b30, 32'h42562399} /* (26, 9, 6) {real, imag} */,
  {32'hc011dd30, 32'h3c2a8000} /* (26, 9, 5) {real, imag} */,
  {32'h42c252f7, 32'h428ba487} /* (26, 9, 4) {real, imag} */,
  {32'h423f8efe, 32'h42bc90ac} /* (26, 9, 3) {real, imag} */,
  {32'hc349e8c3, 32'hc2e3576b} /* (26, 9, 2) {real, imag} */,
  {32'h4200fae0, 32'hc3aaa79f} /* (26, 9, 1) {real, imag} */,
  {32'hc401093c, 32'h00000000} /* (26, 9, 0) {real, imag} */,
  {32'hc2abcfac, 32'h4401c748} /* (26, 8, 31) {real, imag} */,
  {32'hc376ee8d, 32'h43311949} /* (26, 8, 30) {real, imag} */,
  {32'h4250c221, 32'hc2cf261e} /* (26, 8, 29) {real, imag} */,
  {32'h4285aa46, 32'hc25e7933} /* (26, 8, 28) {real, imag} */,
  {32'hc24a18b4, 32'h42124384} /* (26, 8, 27) {real, imag} */,
  {32'hc183bebc, 32'hc1eaa482} /* (26, 8, 26) {real, imag} */,
  {32'h4115a348, 32'hc20d4e0e} /* (26, 8, 25) {real, imag} */,
  {32'hc177f294, 32'hc1c68e6d} /* (26, 8, 24) {real, imag} */,
  {32'hc2a91809, 32'hc226cc8f} /* (26, 8, 23) {real, imag} */,
  {32'hc19d0264, 32'h409cf89c} /* (26, 8, 22) {real, imag} */,
  {32'hc289ca2c, 32'h42071e20} /* (26, 8, 21) {real, imag} */,
  {32'hc2a7c8da, 32'h4225c3d2} /* (26, 8, 20) {real, imag} */,
  {32'hc2606a28, 32'hc130add0} /* (26, 8, 19) {real, imag} */,
  {32'hc1cfcf28, 32'hc1ade184} /* (26, 8, 18) {real, imag} */,
  {32'h412e0a4e, 32'hc1420798} /* (26, 8, 17) {real, imag} */,
  {32'hc17df8df, 32'h00000000} /* (26, 8, 16) {real, imag} */,
  {32'h412e0a4e, 32'h41420798} /* (26, 8, 15) {real, imag} */,
  {32'hc1cfcf28, 32'h41ade184} /* (26, 8, 14) {real, imag} */,
  {32'hc2606a28, 32'h4130add0} /* (26, 8, 13) {real, imag} */,
  {32'hc2a7c8da, 32'hc225c3d2} /* (26, 8, 12) {real, imag} */,
  {32'hc289ca2c, 32'hc2071e20} /* (26, 8, 11) {real, imag} */,
  {32'hc19d0264, 32'hc09cf89c} /* (26, 8, 10) {real, imag} */,
  {32'hc2a91809, 32'h4226cc8f} /* (26, 8, 9) {real, imag} */,
  {32'hc177f294, 32'h41c68e6d} /* (26, 8, 8) {real, imag} */,
  {32'h4115a348, 32'h420d4e0e} /* (26, 8, 7) {real, imag} */,
  {32'hc183bebc, 32'h41eaa482} /* (26, 8, 6) {real, imag} */,
  {32'hc24a18b4, 32'hc2124384} /* (26, 8, 5) {real, imag} */,
  {32'h4285aa46, 32'h425e7933} /* (26, 8, 4) {real, imag} */,
  {32'h4250c221, 32'h42cf261e} /* (26, 8, 3) {real, imag} */,
  {32'hc376ee8d, 32'hc3311949} /* (26, 8, 2) {real, imag} */,
  {32'hc2abcfac, 32'hc401c748} /* (26, 8, 1) {real, imag} */,
  {32'hc46d2ab8, 32'h00000000} /* (26, 8, 0) {real, imag} */,
  {32'hc3a98776, 32'h4409d31e} /* (26, 7, 31) {real, imag} */,
  {32'hc3659f94, 32'h436dae10} /* (26, 7, 30) {real, imag} */,
  {32'h42c7dbf1, 32'h429a1000} /* (26, 7, 29) {real, imag} */,
  {32'h4296c414, 32'hc2a13ae3} /* (26, 7, 28) {real, imag} */,
  {32'h42125725, 32'h414647f8} /* (26, 7, 27) {real, imag} */,
  {32'hc162c206, 32'hc2dca0a4} /* (26, 7, 26) {real, imag} */,
  {32'h42cd3855, 32'hc258c8be} /* (26, 7, 25) {real, imag} */,
  {32'hc28cefa4, 32'hc254e7e2} /* (26, 7, 24) {real, imag} */,
  {32'hc2a0b5e8, 32'h4231f6dc} /* (26, 7, 23) {real, imag} */,
  {32'h429c3afb, 32'h429a982c} /* (26, 7, 22) {real, imag} */,
  {32'h4237cc69, 32'h42db8bac} /* (26, 7, 21) {real, imag} */,
  {32'hc25ebb7a, 32'h424fa38a} /* (26, 7, 20) {real, imag} */,
  {32'h41e4621f, 32'hc157fad6} /* (26, 7, 19) {real, imag} */,
  {32'h410a9bb0, 32'h42185c72} /* (26, 7, 18) {real, imag} */,
  {32'h41cb362c, 32'hc144d8fc} /* (26, 7, 17) {real, imag} */,
  {32'h424b656e, 32'h00000000} /* (26, 7, 16) {real, imag} */,
  {32'h41cb362c, 32'h4144d8fc} /* (26, 7, 15) {real, imag} */,
  {32'h410a9bb0, 32'hc2185c72} /* (26, 7, 14) {real, imag} */,
  {32'h41e4621f, 32'h4157fad6} /* (26, 7, 13) {real, imag} */,
  {32'hc25ebb7a, 32'hc24fa38a} /* (26, 7, 12) {real, imag} */,
  {32'h4237cc69, 32'hc2db8bac} /* (26, 7, 11) {real, imag} */,
  {32'h429c3afb, 32'hc29a982c} /* (26, 7, 10) {real, imag} */,
  {32'hc2a0b5e8, 32'hc231f6dc} /* (26, 7, 9) {real, imag} */,
  {32'hc28cefa4, 32'h4254e7e2} /* (26, 7, 8) {real, imag} */,
  {32'h42cd3855, 32'h4258c8be} /* (26, 7, 7) {real, imag} */,
  {32'hc162c206, 32'h42dca0a4} /* (26, 7, 6) {real, imag} */,
  {32'h42125725, 32'hc14647f8} /* (26, 7, 5) {real, imag} */,
  {32'h4296c414, 32'h42a13ae3} /* (26, 7, 4) {real, imag} */,
  {32'h42c7dbf1, 32'hc29a1000} /* (26, 7, 3) {real, imag} */,
  {32'hc3659f94, 32'hc36dae10} /* (26, 7, 2) {real, imag} */,
  {32'hc3a98776, 32'hc409d31e} /* (26, 7, 1) {real, imag} */,
  {32'hc48fb8a1, 32'h00000000} /* (26, 7, 0) {real, imag} */,
  {32'hc406fcf4, 32'h43fe8648} /* (26, 6, 31) {real, imag} */,
  {32'hc3844aa0, 32'h42dce53d} /* (26, 6, 30) {real, imag} */,
  {32'h42714b32, 32'h41c19379} /* (26, 6, 29) {real, imag} */,
  {32'h42923531, 32'h415bd124} /* (26, 6, 28) {real, imag} */,
  {32'hc17984c6, 32'h42883e57} /* (26, 6, 27) {real, imag} */,
  {32'h417556cf, 32'hc2e105b3} /* (26, 6, 26) {real, imag} */,
  {32'h41873b1b, 32'hc2a2b844} /* (26, 6, 25) {real, imag} */,
  {32'hc21cd946, 32'h413c0b24} /* (26, 6, 24) {real, imag} */,
  {32'h425547aa, 32'h42d271eb} /* (26, 6, 23) {real, imag} */,
  {32'h412ac11a, 32'hc24eeece} /* (26, 6, 22) {real, imag} */,
  {32'hc0ab72a0, 32'hc191578f} /* (26, 6, 21) {real, imag} */,
  {32'hc1d51457, 32'hc2a8ecec} /* (26, 6, 20) {real, imag} */,
  {32'h41a9e4c3, 32'hc1f9ea04} /* (26, 6, 19) {real, imag} */,
  {32'h42049486, 32'hc0bacf74} /* (26, 6, 18) {real, imag} */,
  {32'hc21c7ca9, 32'hc2fe7215} /* (26, 6, 17) {real, imag} */,
  {32'h41d24927, 32'h00000000} /* (26, 6, 16) {real, imag} */,
  {32'hc21c7ca9, 32'h42fe7215} /* (26, 6, 15) {real, imag} */,
  {32'h42049486, 32'h40bacf74} /* (26, 6, 14) {real, imag} */,
  {32'h41a9e4c3, 32'h41f9ea04} /* (26, 6, 13) {real, imag} */,
  {32'hc1d51457, 32'h42a8ecec} /* (26, 6, 12) {real, imag} */,
  {32'hc0ab72a0, 32'h4191578f} /* (26, 6, 11) {real, imag} */,
  {32'h412ac11a, 32'h424eeece} /* (26, 6, 10) {real, imag} */,
  {32'h425547aa, 32'hc2d271eb} /* (26, 6, 9) {real, imag} */,
  {32'hc21cd946, 32'hc13c0b24} /* (26, 6, 8) {real, imag} */,
  {32'h41873b1b, 32'h42a2b844} /* (26, 6, 7) {real, imag} */,
  {32'h417556cf, 32'h42e105b3} /* (26, 6, 6) {real, imag} */,
  {32'hc17984c6, 32'hc2883e57} /* (26, 6, 5) {real, imag} */,
  {32'h42923531, 32'hc15bd124} /* (26, 6, 4) {real, imag} */,
  {32'h42714b32, 32'hc1c19379} /* (26, 6, 3) {real, imag} */,
  {32'hc3844aa0, 32'hc2dce53d} /* (26, 6, 2) {real, imag} */,
  {32'hc406fcf4, 32'hc3fe8648} /* (26, 6, 1) {real, imag} */,
  {32'hc4948b00, 32'h00000000} /* (26, 6, 0) {real, imag} */,
  {32'hc420634e, 32'h4402ab2d} /* (26, 5, 31) {real, imag} */,
  {32'hc2f8fb91, 32'h43136828} /* (26, 5, 30) {real, imag} */,
  {32'h430ff71e, 32'hc3088b26} /* (26, 5, 29) {real, imag} */,
  {32'h4220c722, 32'h42a4ebf1} /* (26, 5, 28) {real, imag} */,
  {32'hc2a5037e, 32'h432c4082} /* (26, 5, 27) {real, imag} */,
  {32'h410258c0, 32'h4185bc6c} /* (26, 5, 26) {real, imag} */,
  {32'h4209da75, 32'hc16cae28} /* (26, 5, 25) {real, imag} */,
  {32'h42c26dbe, 32'h42d9d210} /* (26, 5, 24) {real, imag} */,
  {32'h4152843a, 32'h4161a4ec} /* (26, 5, 23) {real, imag} */,
  {32'hc1a57394, 32'h429bae3a} /* (26, 5, 22) {real, imag} */,
  {32'h427653f5, 32'h41c84eba} /* (26, 5, 21) {real, imag} */,
  {32'hc0dc7ed8, 32'h41eab128} /* (26, 5, 20) {real, imag} */,
  {32'hbe3c3000, 32'hc2aa9d3a} /* (26, 5, 19) {real, imag} */,
  {32'hc1833c36, 32'h4325c61a} /* (26, 5, 18) {real, imag} */,
  {32'hc20b0263, 32'hc17b19a8} /* (26, 5, 17) {real, imag} */,
  {32'hc2cb8734, 32'h00000000} /* (26, 5, 16) {real, imag} */,
  {32'hc20b0263, 32'h417b19a8} /* (26, 5, 15) {real, imag} */,
  {32'hc1833c36, 32'hc325c61a} /* (26, 5, 14) {real, imag} */,
  {32'hbe3c3000, 32'h42aa9d3a} /* (26, 5, 13) {real, imag} */,
  {32'hc0dc7ed8, 32'hc1eab128} /* (26, 5, 12) {real, imag} */,
  {32'h427653f5, 32'hc1c84eba} /* (26, 5, 11) {real, imag} */,
  {32'hc1a57394, 32'hc29bae3a} /* (26, 5, 10) {real, imag} */,
  {32'h4152843a, 32'hc161a4ec} /* (26, 5, 9) {real, imag} */,
  {32'h42c26dbe, 32'hc2d9d210} /* (26, 5, 8) {real, imag} */,
  {32'h4209da75, 32'h416cae28} /* (26, 5, 7) {real, imag} */,
  {32'h410258c0, 32'hc185bc6c} /* (26, 5, 6) {real, imag} */,
  {32'hc2a5037e, 32'hc32c4082} /* (26, 5, 5) {real, imag} */,
  {32'h4220c722, 32'hc2a4ebf1} /* (26, 5, 4) {real, imag} */,
  {32'h430ff71e, 32'h43088b26} /* (26, 5, 3) {real, imag} */,
  {32'hc2f8fb91, 32'hc3136828} /* (26, 5, 2) {real, imag} */,
  {32'hc420634e, 32'hc402ab2d} /* (26, 5, 1) {real, imag} */,
  {32'hc4b7875f, 32'h00000000} /* (26, 5, 0) {real, imag} */,
  {32'hc4453b70, 32'h4428806b} /* (26, 4, 31) {real, imag} */,
  {32'hc20196be, 32'h438460fe} /* (26, 4, 30) {real, imag} */,
  {32'h4287c1ec, 32'h423c265e} /* (26, 4, 29) {real, imag} */,
  {32'hc2abab9c, 32'hc209e314} /* (26, 4, 28) {real, imag} */,
  {32'hc21c5d3d, 32'h42850e7c} /* (26, 4, 27) {real, imag} */,
  {32'h430eea84, 32'hc242b306} /* (26, 4, 26) {real, imag} */,
  {32'hc29ced9c, 32'hc2b3a374} /* (26, 4, 25) {real, imag} */,
  {32'h42240274, 32'h42c33eed} /* (26, 4, 24) {real, imag} */,
  {32'hbfc5ace8, 32'h42d34df6} /* (26, 4, 23) {real, imag} */,
  {32'hc272724a, 32'h4173fac0} /* (26, 4, 22) {real, imag} */,
  {32'hc28df848, 32'h40322fe5} /* (26, 4, 21) {real, imag} */,
  {32'h42524acc, 32'hc3254b95} /* (26, 4, 20) {real, imag} */,
  {32'h41a505f0, 32'h41c12d52} /* (26, 4, 19) {real, imag} */,
  {32'h40c3e42c, 32'hc129f3d4} /* (26, 4, 18) {real, imag} */,
  {32'h422f7a91, 32'h4137d8f6} /* (26, 4, 17) {real, imag} */,
  {32'hc14b6144, 32'h00000000} /* (26, 4, 16) {real, imag} */,
  {32'h422f7a91, 32'hc137d8f6} /* (26, 4, 15) {real, imag} */,
  {32'h40c3e42c, 32'h4129f3d4} /* (26, 4, 14) {real, imag} */,
  {32'h41a505f0, 32'hc1c12d52} /* (26, 4, 13) {real, imag} */,
  {32'h42524acc, 32'h43254b95} /* (26, 4, 12) {real, imag} */,
  {32'hc28df848, 32'hc0322fe5} /* (26, 4, 11) {real, imag} */,
  {32'hc272724a, 32'hc173fac0} /* (26, 4, 10) {real, imag} */,
  {32'hbfc5ace8, 32'hc2d34df6} /* (26, 4, 9) {real, imag} */,
  {32'h42240274, 32'hc2c33eed} /* (26, 4, 8) {real, imag} */,
  {32'hc29ced9c, 32'h42b3a374} /* (26, 4, 7) {real, imag} */,
  {32'h430eea84, 32'h4242b306} /* (26, 4, 6) {real, imag} */,
  {32'hc21c5d3d, 32'hc2850e7c} /* (26, 4, 5) {real, imag} */,
  {32'hc2abab9c, 32'h4209e314} /* (26, 4, 4) {real, imag} */,
  {32'h4287c1ec, 32'hc23c265e} /* (26, 4, 3) {real, imag} */,
  {32'hc20196be, 32'hc38460fe} /* (26, 4, 2) {real, imag} */,
  {32'hc4453b70, 32'hc428806b} /* (26, 4, 1) {real, imag} */,
  {32'hc4ac1a02, 32'h00000000} /* (26, 4, 0) {real, imag} */,
  {32'hc451b1e5, 32'h4433b479} /* (26, 3, 31) {real, imag} */,
  {32'h42cca584, 32'h4389e80b} /* (26, 3, 30) {real, imag} */,
  {32'hc148e8c4, 32'hc12b4b88} /* (26, 3, 29) {real, imag} */,
  {32'hc240de5f, 32'h41397ae4} /* (26, 3, 28) {real, imag} */,
  {32'h4166db30, 32'hc1814e76} /* (26, 3, 27) {real, imag} */,
  {32'h41d64fee, 32'h41e23344} /* (26, 3, 26) {real, imag} */,
  {32'hc2f59ab1, 32'hc1dbb31d} /* (26, 3, 25) {real, imag} */,
  {32'hc29e49ac, 32'hc2ccbdf4} /* (26, 3, 24) {real, imag} */,
  {32'h41d74170, 32'h431aa435} /* (26, 3, 23) {real, imag} */,
  {32'hc3039220, 32'hc2662e24} /* (26, 3, 22) {real, imag} */,
  {32'hc2dfd85a, 32'hc1dc4d6c} /* (26, 3, 21) {real, imag} */,
  {32'h4117a788, 32'hc144a482} /* (26, 3, 20) {real, imag} */,
  {32'h4245855f, 32'h42223db2} /* (26, 3, 19) {real, imag} */,
  {32'h42efa126, 32'h4186b054} /* (26, 3, 18) {real, imag} */,
  {32'h409c9650, 32'h430c8bea} /* (26, 3, 17) {real, imag} */,
  {32'h42ae06d8, 32'h00000000} /* (26, 3, 16) {real, imag} */,
  {32'h409c9650, 32'hc30c8bea} /* (26, 3, 15) {real, imag} */,
  {32'h42efa126, 32'hc186b054} /* (26, 3, 14) {real, imag} */,
  {32'h4245855f, 32'hc2223db2} /* (26, 3, 13) {real, imag} */,
  {32'h4117a788, 32'h4144a482} /* (26, 3, 12) {real, imag} */,
  {32'hc2dfd85a, 32'h41dc4d6c} /* (26, 3, 11) {real, imag} */,
  {32'hc3039220, 32'h42662e24} /* (26, 3, 10) {real, imag} */,
  {32'h41d74170, 32'hc31aa435} /* (26, 3, 9) {real, imag} */,
  {32'hc29e49ac, 32'h42ccbdf4} /* (26, 3, 8) {real, imag} */,
  {32'hc2f59ab1, 32'h41dbb31d} /* (26, 3, 7) {real, imag} */,
  {32'h41d64fee, 32'hc1e23344} /* (26, 3, 6) {real, imag} */,
  {32'h4166db30, 32'h41814e76} /* (26, 3, 5) {real, imag} */,
  {32'hc240de5f, 32'hc1397ae4} /* (26, 3, 4) {real, imag} */,
  {32'hc148e8c4, 32'h412b4b88} /* (26, 3, 3) {real, imag} */,
  {32'h42cca584, 32'hc389e80b} /* (26, 3, 2) {real, imag} */,
  {32'hc451b1e5, 32'hc433b479} /* (26, 3, 1) {real, imag} */,
  {32'hc4a6cb3b, 32'h00000000} /* (26, 3, 0) {real, imag} */,
  {32'hc46b0f8b, 32'h43f7262d} /* (26, 2, 31) {real, imag} */,
  {32'h4348914e, 32'h4344d468} /* (26, 2, 30) {real, imag} */,
  {32'h41e359d0, 32'hc0d90814} /* (26, 2, 29) {real, imag} */,
  {32'h430ba30b, 32'hbfc6c5b8} /* (26, 2, 28) {real, imag} */,
  {32'hc29848bc, 32'hc19e13f4} /* (26, 2, 27) {real, imag} */,
  {32'hc280b7a6, 32'hc24bd1fe} /* (26, 2, 26) {real, imag} */,
  {32'hc2d15d78, 32'hc2008d62} /* (26, 2, 25) {real, imag} */,
  {32'hc2801892, 32'h4125889c} /* (26, 2, 24) {real, imag} */,
  {32'hc1599ffc, 32'hc2aa6742} /* (26, 2, 23) {real, imag} */,
  {32'hc1434317, 32'h41ed0608} /* (26, 2, 22) {real, imag} */,
  {32'hc0a1d950, 32'h42b1237e} /* (26, 2, 21) {real, imag} */,
  {32'hc1d9ade5, 32'h402cb040} /* (26, 2, 20) {real, imag} */,
  {32'h4208cc42, 32'hc26dec86} /* (26, 2, 19) {real, imag} */,
  {32'h41b428b6, 32'h427b3b94} /* (26, 2, 18) {real, imag} */,
  {32'h42364a60, 32'h4152296e} /* (26, 2, 17) {real, imag} */,
  {32'hc1b8ba92, 32'h00000000} /* (26, 2, 16) {real, imag} */,
  {32'h42364a60, 32'hc152296e} /* (26, 2, 15) {real, imag} */,
  {32'h41b428b6, 32'hc27b3b94} /* (26, 2, 14) {real, imag} */,
  {32'h4208cc42, 32'h426dec86} /* (26, 2, 13) {real, imag} */,
  {32'hc1d9ade5, 32'hc02cb040} /* (26, 2, 12) {real, imag} */,
  {32'hc0a1d950, 32'hc2b1237e} /* (26, 2, 11) {real, imag} */,
  {32'hc1434317, 32'hc1ed0608} /* (26, 2, 10) {real, imag} */,
  {32'hc1599ffc, 32'h42aa6742} /* (26, 2, 9) {real, imag} */,
  {32'hc2801892, 32'hc125889c} /* (26, 2, 8) {real, imag} */,
  {32'hc2d15d78, 32'h42008d62} /* (26, 2, 7) {real, imag} */,
  {32'hc280b7a6, 32'h424bd1fe} /* (26, 2, 6) {real, imag} */,
  {32'hc29848bc, 32'h419e13f4} /* (26, 2, 5) {real, imag} */,
  {32'h430ba30b, 32'h3fc6c5b8} /* (26, 2, 4) {real, imag} */,
  {32'h41e359d0, 32'h40d90814} /* (26, 2, 3) {real, imag} */,
  {32'h4348914e, 32'hc344d468} /* (26, 2, 2) {real, imag} */,
  {32'hc46b0f8b, 32'hc3f7262d} /* (26, 2, 1) {real, imag} */,
  {32'hc4b5f61c, 32'h00000000} /* (26, 2, 0) {real, imag} */,
  {32'hc46deb28, 32'h43d6de96} /* (26, 1, 31) {real, imag} */,
  {32'h42e81329, 32'h434af277} /* (26, 1, 30) {real, imag} */,
  {32'hc1992480, 32'h4281191a} /* (26, 1, 29) {real, imag} */,
  {32'h414d908a, 32'h4323eef5} /* (26, 1, 28) {real, imag} */,
  {32'hc2599990, 32'hc2fa2f03} /* (26, 1, 27) {real, imag} */,
  {32'hc2997bfe, 32'hc1e4808e} /* (26, 1, 26) {real, imag} */,
  {32'hc2aa9ebf, 32'hc309fea2} /* (26, 1, 25) {real, imag} */,
  {32'h43215784, 32'hc1f09c74} /* (26, 1, 24) {real, imag} */,
  {32'hc231afc7, 32'hc1358602} /* (26, 1, 23) {real, imag} */,
  {32'hc219a3d0, 32'h430c8458} /* (26, 1, 22) {real, imag} */,
  {32'hc2227382, 32'hc2230f88} /* (26, 1, 21) {real, imag} */,
  {32'h41c5ae84, 32'h4216be76} /* (26, 1, 20) {real, imag} */,
  {32'h4247c1d8, 32'hc25adef9} /* (26, 1, 19) {real, imag} */,
  {32'hc15dde2a, 32'hc26d5665} /* (26, 1, 18) {real, imag} */,
  {32'h41b34e8e, 32'h421e6c20} /* (26, 1, 17) {real, imag} */,
  {32'h416faf30, 32'h00000000} /* (26, 1, 16) {real, imag} */,
  {32'h41b34e8e, 32'hc21e6c20} /* (26, 1, 15) {real, imag} */,
  {32'hc15dde2a, 32'h426d5665} /* (26, 1, 14) {real, imag} */,
  {32'h4247c1d8, 32'h425adef9} /* (26, 1, 13) {real, imag} */,
  {32'h41c5ae84, 32'hc216be76} /* (26, 1, 12) {real, imag} */,
  {32'hc2227382, 32'h42230f88} /* (26, 1, 11) {real, imag} */,
  {32'hc219a3d0, 32'hc30c8458} /* (26, 1, 10) {real, imag} */,
  {32'hc231afc7, 32'h41358602} /* (26, 1, 9) {real, imag} */,
  {32'h43215784, 32'h41f09c74} /* (26, 1, 8) {real, imag} */,
  {32'hc2aa9ebf, 32'h4309fea2} /* (26, 1, 7) {real, imag} */,
  {32'hc2997bfe, 32'h41e4808e} /* (26, 1, 6) {real, imag} */,
  {32'hc2599990, 32'h42fa2f03} /* (26, 1, 5) {real, imag} */,
  {32'h414d908a, 32'hc323eef5} /* (26, 1, 4) {real, imag} */,
  {32'hc1992480, 32'hc281191a} /* (26, 1, 3) {real, imag} */,
  {32'h42e81329, 32'hc34af277} /* (26, 1, 2) {real, imag} */,
  {32'hc46deb28, 32'hc3d6de96} /* (26, 1, 1) {real, imag} */,
  {32'hc4cb48ff, 32'h00000000} /* (26, 1, 0) {real, imag} */,
  {32'hc4818b32, 32'h43c2ade1} /* (26, 0, 31) {real, imag} */,
  {32'h431332fc, 32'h43626c02} /* (26, 0, 30) {real, imag} */,
  {32'h424fde4c, 32'hc2857d43} /* (26, 0, 29) {real, imag} */,
  {32'hc289d1f7, 32'h42b986e7} /* (26, 0, 28) {real, imag} */,
  {32'hbf8fc5a0, 32'hc29e6e62} /* (26, 0, 27) {real, imag} */,
  {32'hc2876c0e, 32'hc297980d} /* (26, 0, 26) {real, imag} */,
  {32'h424d1946, 32'hc20d00d8} /* (26, 0, 25) {real, imag} */,
  {32'h4251f71b, 32'h4158d362} /* (26, 0, 24) {real, imag} */,
  {32'hc1c3f209, 32'h4259215b} /* (26, 0, 23) {real, imag} */,
  {32'hc25dd3f8, 32'h429a9ae4} /* (26, 0, 22) {real, imag} */,
  {32'h42865a02, 32'hc2c12f73} /* (26, 0, 21) {real, imag} */,
  {32'hc178b6da, 32'h424b0150} /* (26, 0, 20) {real, imag} */,
  {32'h41b0a887, 32'h424bdd1e} /* (26, 0, 19) {real, imag} */,
  {32'hc18afd8e, 32'hc1d80ab8} /* (26, 0, 18) {real, imag} */,
  {32'h41fe97e0, 32'h41031bea} /* (26, 0, 17) {real, imag} */,
  {32'h420b125b, 32'h00000000} /* (26, 0, 16) {real, imag} */,
  {32'h41fe97e0, 32'hc1031bea} /* (26, 0, 15) {real, imag} */,
  {32'hc18afd8e, 32'h41d80ab8} /* (26, 0, 14) {real, imag} */,
  {32'h41b0a887, 32'hc24bdd1e} /* (26, 0, 13) {real, imag} */,
  {32'hc178b6da, 32'hc24b0150} /* (26, 0, 12) {real, imag} */,
  {32'h42865a02, 32'h42c12f73} /* (26, 0, 11) {real, imag} */,
  {32'hc25dd3f8, 32'hc29a9ae4} /* (26, 0, 10) {real, imag} */,
  {32'hc1c3f209, 32'hc259215b} /* (26, 0, 9) {real, imag} */,
  {32'h4251f71b, 32'hc158d362} /* (26, 0, 8) {real, imag} */,
  {32'h424d1946, 32'h420d00d8} /* (26, 0, 7) {real, imag} */,
  {32'hc2876c0e, 32'h4297980d} /* (26, 0, 6) {real, imag} */,
  {32'hbf8fc5a0, 32'h429e6e62} /* (26, 0, 5) {real, imag} */,
  {32'hc289d1f7, 32'hc2b986e7} /* (26, 0, 4) {real, imag} */,
  {32'h424fde4c, 32'h42857d43} /* (26, 0, 3) {real, imag} */,
  {32'h431332fc, 32'hc3626c02} /* (26, 0, 2) {real, imag} */,
  {32'hc4818b32, 32'hc3c2ade1} /* (26, 0, 1) {real, imag} */,
  {32'hc4dc00a2, 32'h00000000} /* (26, 0, 0) {real, imag} */,
  {32'hc50961c9, 32'h448b1db2} /* (25, 31, 31) {real, imag} */,
  {32'h43b05348, 32'hc2a757a0} /* (25, 31, 30) {real, imag} */,
  {32'h41c54dc8, 32'hc261b76c} /* (25, 31, 29) {real, imag} */,
  {32'hc2cc5927, 32'h4220f477} /* (25, 31, 28) {real, imag} */,
  {32'h42f5693e, 32'hc2535b12} /* (25, 31, 27) {real, imag} */,
  {32'hc23c1afd, 32'hc1ee7101} /* (25, 31, 26) {real, imag} */,
  {32'h41bc4d13, 32'hc2008fc7} /* (25, 31, 25) {real, imag} */,
  {32'hc1b42420, 32'hc20a042c} /* (25, 31, 24) {real, imag} */,
  {32'hc140000e, 32'hc26faca2} /* (25, 31, 23) {real, imag} */,
  {32'h41900c16, 32'hc20f15b0} /* (25, 31, 22) {real, imag} */,
  {32'h41cebb23, 32'hc1a33f70} /* (25, 31, 21) {real, imag} */,
  {32'h42106217, 32'hc228ffd8} /* (25, 31, 20) {real, imag} */,
  {32'h41899754, 32'hc1810e68} /* (25, 31, 19) {real, imag} */,
  {32'hc2198a7e, 32'hc29eab15} /* (25, 31, 18) {real, imag} */,
  {32'h4235d1ab, 32'hc0febde1} /* (25, 31, 17) {real, imag} */,
  {32'h42900102, 32'h00000000} /* (25, 31, 16) {real, imag} */,
  {32'h4235d1ab, 32'h40febde1} /* (25, 31, 15) {real, imag} */,
  {32'hc2198a7e, 32'h429eab15} /* (25, 31, 14) {real, imag} */,
  {32'h41899754, 32'h41810e68} /* (25, 31, 13) {real, imag} */,
  {32'h42106217, 32'h4228ffd8} /* (25, 31, 12) {real, imag} */,
  {32'h41cebb23, 32'h41a33f70} /* (25, 31, 11) {real, imag} */,
  {32'h41900c16, 32'h420f15b0} /* (25, 31, 10) {real, imag} */,
  {32'hc140000e, 32'h426faca2} /* (25, 31, 9) {real, imag} */,
  {32'hc1b42420, 32'h420a042c} /* (25, 31, 8) {real, imag} */,
  {32'h41bc4d13, 32'h42008fc7} /* (25, 31, 7) {real, imag} */,
  {32'hc23c1afd, 32'h41ee7101} /* (25, 31, 6) {real, imag} */,
  {32'h42f5693e, 32'h42535b12} /* (25, 31, 5) {real, imag} */,
  {32'hc2cc5927, 32'hc220f477} /* (25, 31, 4) {real, imag} */,
  {32'h41c54dc8, 32'h4261b76c} /* (25, 31, 3) {real, imag} */,
  {32'h43b05348, 32'h42a757a0} /* (25, 31, 2) {real, imag} */,
  {32'hc50961c9, 32'hc48b1db2} /* (25, 31, 1) {real, imag} */,
  {32'hc542c599, 32'h00000000} /* (25, 31, 0) {real, imag} */,
  {32'hc51d84de, 32'h4473df27} /* (25, 30, 31) {real, imag} */,
  {32'h442a8dc4, 32'hc2bdb9de} /* (25, 30, 30) {real, imag} */,
  {32'h412ec19c, 32'hc29e42a6} /* (25, 30, 29) {real, imag} */,
  {32'hc31b58ea, 32'h42132898} /* (25, 30, 28) {real, imag} */,
  {32'h42b9cd31, 32'h419dde35} /* (25, 30, 27) {real, imag} */,
  {32'h422ac3b1, 32'hc26db6d0} /* (25, 30, 26) {real, imag} */,
  {32'hc1887d86, 32'hc28575be} /* (25, 30, 25) {real, imag} */,
  {32'hc0aa9000, 32'hc2233490} /* (25, 30, 24) {real, imag} */,
  {32'hc214a523, 32'hc1c27966} /* (25, 30, 23) {real, imag} */,
  {32'hc135aab0, 32'hc235ea96} /* (25, 30, 22) {real, imag} */,
  {32'hc22d3a9b, 32'hc202a03a} /* (25, 30, 21) {real, imag} */,
  {32'h41bf991d, 32'hc2074dca} /* (25, 30, 20) {real, imag} */,
  {32'h426eac27, 32'h426fbabe} /* (25, 30, 19) {real, imag} */,
  {32'h41cc18cc, 32'hc2f098ec} /* (25, 30, 18) {real, imag} */,
  {32'hc104d3ca, 32'h41937209} /* (25, 30, 17) {real, imag} */,
  {32'hc0db080c, 32'h00000000} /* (25, 30, 16) {real, imag} */,
  {32'hc104d3ca, 32'hc1937209} /* (25, 30, 15) {real, imag} */,
  {32'h41cc18cc, 32'h42f098ec} /* (25, 30, 14) {real, imag} */,
  {32'h426eac27, 32'hc26fbabe} /* (25, 30, 13) {real, imag} */,
  {32'h41bf991d, 32'h42074dca} /* (25, 30, 12) {real, imag} */,
  {32'hc22d3a9b, 32'h4202a03a} /* (25, 30, 11) {real, imag} */,
  {32'hc135aab0, 32'h4235ea96} /* (25, 30, 10) {real, imag} */,
  {32'hc214a523, 32'h41c27966} /* (25, 30, 9) {real, imag} */,
  {32'hc0aa9000, 32'h42233490} /* (25, 30, 8) {real, imag} */,
  {32'hc1887d86, 32'h428575be} /* (25, 30, 7) {real, imag} */,
  {32'h422ac3b1, 32'h426db6d0} /* (25, 30, 6) {real, imag} */,
  {32'h42b9cd31, 32'hc19dde35} /* (25, 30, 5) {real, imag} */,
  {32'hc31b58ea, 32'hc2132898} /* (25, 30, 4) {real, imag} */,
  {32'h412ec19c, 32'h429e42a6} /* (25, 30, 3) {real, imag} */,
  {32'h442a8dc4, 32'h42bdb9de} /* (25, 30, 2) {real, imag} */,
  {32'hc51d84de, 32'hc473df27} /* (25, 30, 1) {real, imag} */,
  {32'hc546139e, 32'h00000000} /* (25, 30, 0) {real, imag} */,
  {32'hc5189312, 32'h4478aeba} /* (25, 29, 31) {real, imag} */,
  {32'h4437246a, 32'h41ddd080} /* (25, 29, 30) {real, imag} */,
  {32'h420db360, 32'hc299bbf2} /* (25, 29, 29) {real, imag} */,
  {32'hc31202fb, 32'hc22b796e} /* (25, 29, 28) {real, imag} */,
  {32'h4299ba3a, 32'hc3560870} /* (25, 29, 27) {real, imag} */,
  {32'h421907de, 32'hc16bbe30} /* (25, 29, 26) {real, imag} */,
  {32'h4323807c, 32'h42ec21fc} /* (25, 29, 25) {real, imag} */,
  {32'h430185f6, 32'hc20f8b82} /* (25, 29, 24) {real, imag} */,
  {32'h40c90a28, 32'h41f05e3a} /* (25, 29, 23) {real, imag} */,
  {32'hc1632fc0, 32'h41319ab6} /* (25, 29, 22) {real, imag} */,
  {32'h42cf4648, 32'hc2bb9e20} /* (25, 29, 21) {real, imag} */,
  {32'hc2b4e1d3, 32'h429336f3} /* (25, 29, 20) {real, imag} */,
  {32'h415cde76, 32'h42166031} /* (25, 29, 19) {real, imag} */,
  {32'h4189b7ec, 32'hc2945c67} /* (25, 29, 18) {real, imag} */,
  {32'hc049d898, 32'h4249428c} /* (25, 29, 17) {real, imag} */,
  {32'h41aaf559, 32'h00000000} /* (25, 29, 16) {real, imag} */,
  {32'hc049d898, 32'hc249428c} /* (25, 29, 15) {real, imag} */,
  {32'h4189b7ec, 32'h42945c67} /* (25, 29, 14) {real, imag} */,
  {32'h415cde76, 32'hc2166031} /* (25, 29, 13) {real, imag} */,
  {32'hc2b4e1d3, 32'hc29336f3} /* (25, 29, 12) {real, imag} */,
  {32'h42cf4648, 32'h42bb9e20} /* (25, 29, 11) {real, imag} */,
  {32'hc1632fc0, 32'hc1319ab6} /* (25, 29, 10) {real, imag} */,
  {32'h40c90a28, 32'hc1f05e3a} /* (25, 29, 9) {real, imag} */,
  {32'h430185f6, 32'h420f8b82} /* (25, 29, 8) {real, imag} */,
  {32'h4323807c, 32'hc2ec21fc} /* (25, 29, 7) {real, imag} */,
  {32'h421907de, 32'h416bbe30} /* (25, 29, 6) {real, imag} */,
  {32'h4299ba3a, 32'h43560870} /* (25, 29, 5) {real, imag} */,
  {32'hc31202fb, 32'h422b796e} /* (25, 29, 4) {real, imag} */,
  {32'h420db360, 32'h4299bbf2} /* (25, 29, 3) {real, imag} */,
  {32'h4437246a, 32'hc1ddd080} /* (25, 29, 2) {real, imag} */,
  {32'hc5189312, 32'hc478aeba} /* (25, 29, 1) {real, imag} */,
  {32'hc552ed26, 32'h00000000} /* (25, 29, 0) {real, imag} */,
  {32'hc5245522, 32'h44645b0f} /* (25, 28, 31) {real, imag} */,
  {32'h443d98c8, 32'hc24ea7f4} /* (25, 28, 30) {real, imag} */,
  {32'h4173c2f8, 32'hc30a01ee} /* (25, 28, 29) {real, imag} */,
  {32'hc2c21e86, 32'h42d328d6} /* (25, 28, 28) {real, imag} */,
  {32'h42eda673, 32'hc362e26b} /* (25, 28, 27) {real, imag} */,
  {32'hc243ce17, 32'h42d27aac} /* (25, 28, 26) {real, imag} */,
  {32'h427ec37d, 32'h3d2ef100} /* (25, 28, 25) {real, imag} */,
  {32'h41bae4e5, 32'hc305f23d} /* (25, 28, 24) {real, imag} */,
  {32'h42852fa4, 32'hc20d159e} /* (25, 28, 23) {real, imag} */,
  {32'hc0c50308, 32'hc28e2308} /* (25, 28, 22) {real, imag} */,
  {32'h42be1c9d, 32'hc26d9291} /* (25, 28, 21) {real, imag} */,
  {32'hc2b7dcce, 32'hc13ab70e} /* (25, 28, 20) {real, imag} */,
  {32'hc2076798, 32'hc23d0aff} /* (25, 28, 19) {real, imag} */,
  {32'hc19faa06, 32'hc2b3c804} /* (25, 28, 18) {real, imag} */,
  {32'hc28bf7de, 32'h42420dae} /* (25, 28, 17) {real, imag} */,
  {32'h431078eb, 32'h00000000} /* (25, 28, 16) {real, imag} */,
  {32'hc28bf7de, 32'hc2420dae} /* (25, 28, 15) {real, imag} */,
  {32'hc19faa06, 32'h42b3c804} /* (25, 28, 14) {real, imag} */,
  {32'hc2076798, 32'h423d0aff} /* (25, 28, 13) {real, imag} */,
  {32'hc2b7dcce, 32'h413ab70e} /* (25, 28, 12) {real, imag} */,
  {32'h42be1c9d, 32'h426d9291} /* (25, 28, 11) {real, imag} */,
  {32'hc0c50308, 32'h428e2308} /* (25, 28, 10) {real, imag} */,
  {32'h42852fa4, 32'h420d159e} /* (25, 28, 9) {real, imag} */,
  {32'h41bae4e5, 32'h4305f23d} /* (25, 28, 8) {real, imag} */,
  {32'h427ec37d, 32'hbd2ef100} /* (25, 28, 7) {real, imag} */,
  {32'hc243ce17, 32'hc2d27aac} /* (25, 28, 6) {real, imag} */,
  {32'h42eda673, 32'h4362e26b} /* (25, 28, 5) {real, imag} */,
  {32'hc2c21e86, 32'hc2d328d6} /* (25, 28, 4) {real, imag} */,
  {32'h4173c2f8, 32'h430a01ee} /* (25, 28, 3) {real, imag} */,
  {32'h443d98c8, 32'h424ea7f4} /* (25, 28, 2) {real, imag} */,
  {32'hc5245522, 32'hc4645b0f} /* (25, 28, 1) {real, imag} */,
  {32'hc55d778a, 32'h00000000} /* (25, 28, 0) {real, imag} */,
  {32'hc524652c, 32'h4429e4be} /* (25, 27, 31) {real, imag} */,
  {32'h4460413c, 32'hc20be5a0} /* (25, 27, 30) {real, imag} */,
  {32'h4288f712, 32'hc35aade8} /* (25, 27, 29) {real, imag} */,
  {32'hc199afac, 32'hc1f0de7a} /* (25, 27, 28) {real, imag} */,
  {32'h4320e3ea, 32'hc35ec030} /* (25, 27, 27) {real, imag} */,
  {32'h41841904, 32'h431bfa24} /* (25, 27, 26) {real, imag} */,
  {32'hc2655a32, 32'h42d606f3} /* (25, 27, 25) {real, imag} */,
  {32'hc18f89aa, 32'hc30c3170} /* (25, 27, 24) {real, imag} */,
  {32'hc088f9b8, 32'h42802dde} /* (25, 27, 23) {real, imag} */,
  {32'hc205d6ba, 32'h4229069b} /* (25, 27, 22) {real, imag} */,
  {32'hc2560db1, 32'hc2ceabd9} /* (25, 27, 21) {real, imag} */,
  {32'hc1722bc2, 32'hc305ea78} /* (25, 27, 20) {real, imag} */,
  {32'h40ae075a, 32'h42829cc7} /* (25, 27, 19) {real, imag} */,
  {32'hc1b6d184, 32'hc24de5c3} /* (25, 27, 18) {real, imag} */,
  {32'h4125d6cc, 32'hc1784d28} /* (25, 27, 17) {real, imag} */,
  {32'h41741fbc, 32'h00000000} /* (25, 27, 16) {real, imag} */,
  {32'h4125d6cc, 32'h41784d28} /* (25, 27, 15) {real, imag} */,
  {32'hc1b6d184, 32'h424de5c3} /* (25, 27, 14) {real, imag} */,
  {32'h40ae075a, 32'hc2829cc7} /* (25, 27, 13) {real, imag} */,
  {32'hc1722bc2, 32'h4305ea78} /* (25, 27, 12) {real, imag} */,
  {32'hc2560db1, 32'h42ceabd9} /* (25, 27, 11) {real, imag} */,
  {32'hc205d6ba, 32'hc229069b} /* (25, 27, 10) {real, imag} */,
  {32'hc088f9b8, 32'hc2802dde} /* (25, 27, 9) {real, imag} */,
  {32'hc18f89aa, 32'h430c3170} /* (25, 27, 8) {real, imag} */,
  {32'hc2655a32, 32'hc2d606f3} /* (25, 27, 7) {real, imag} */,
  {32'h41841904, 32'hc31bfa24} /* (25, 27, 6) {real, imag} */,
  {32'h4320e3ea, 32'h435ec030} /* (25, 27, 5) {real, imag} */,
  {32'hc199afac, 32'h41f0de7a} /* (25, 27, 4) {real, imag} */,
  {32'h4288f712, 32'h435aade8} /* (25, 27, 3) {real, imag} */,
  {32'h4460413c, 32'h420be5a0} /* (25, 27, 2) {real, imag} */,
  {32'hc524652c, 32'hc429e4be} /* (25, 27, 1) {real, imag} */,
  {32'hc55cb2b2, 32'h00000000} /* (25, 27, 0) {real, imag} */,
  {32'hc51c5f65, 32'h441056ec} /* (25, 26, 31) {real, imag} */,
  {32'h444332d5, 32'h42fb15a9} /* (25, 26, 30) {real, imag} */,
  {32'h419c2794, 32'h41533356} /* (25, 26, 29) {real, imag} */,
  {32'hc1fa292d, 32'h41d61d71} /* (25, 26, 28) {real, imag} */,
  {32'h4305285e, 32'hc318affd} /* (25, 26, 27) {real, imag} */,
  {32'h4253504a, 32'h4231e150} /* (25, 26, 26) {real, imag} */,
  {32'h424f9932, 32'hc090b6f8} /* (25, 26, 25) {real, imag} */,
  {32'hc14b745d, 32'hc34f1450} /* (25, 26, 24) {real, imag} */,
  {32'h3ed23fc0, 32'h40b362d4} /* (25, 26, 23) {real, imag} */,
  {32'h3d55e500, 32'h4246b5d2} /* (25, 26, 22) {real, imag} */,
  {32'hc2023045, 32'h41178c42} /* (25, 26, 21) {real, imag} */,
  {32'h420d7f0c, 32'h41bb44e8} /* (25, 26, 20) {real, imag} */,
  {32'hc2272328, 32'h4200daf8} /* (25, 26, 19) {real, imag} */,
  {32'hc234a3ee, 32'hc1c52eb1} /* (25, 26, 18) {real, imag} */,
  {32'hc19948ec, 32'h40cc3e80} /* (25, 26, 17) {real, imag} */,
  {32'h42cc921b, 32'h00000000} /* (25, 26, 16) {real, imag} */,
  {32'hc19948ec, 32'hc0cc3e80} /* (25, 26, 15) {real, imag} */,
  {32'hc234a3ee, 32'h41c52eb1} /* (25, 26, 14) {real, imag} */,
  {32'hc2272328, 32'hc200daf8} /* (25, 26, 13) {real, imag} */,
  {32'h420d7f0c, 32'hc1bb44e8} /* (25, 26, 12) {real, imag} */,
  {32'hc2023045, 32'hc1178c42} /* (25, 26, 11) {real, imag} */,
  {32'h3d55e500, 32'hc246b5d2} /* (25, 26, 10) {real, imag} */,
  {32'h3ed23fc0, 32'hc0b362d4} /* (25, 26, 9) {real, imag} */,
  {32'hc14b745d, 32'h434f1450} /* (25, 26, 8) {real, imag} */,
  {32'h424f9932, 32'h4090b6f8} /* (25, 26, 7) {real, imag} */,
  {32'h4253504a, 32'hc231e150} /* (25, 26, 6) {real, imag} */,
  {32'h4305285e, 32'h4318affd} /* (25, 26, 5) {real, imag} */,
  {32'hc1fa292d, 32'hc1d61d71} /* (25, 26, 4) {real, imag} */,
  {32'h419c2794, 32'hc1533356} /* (25, 26, 3) {real, imag} */,
  {32'h444332d5, 32'hc2fb15a9} /* (25, 26, 2) {real, imag} */,
  {32'hc51c5f65, 32'hc41056ec} /* (25, 26, 1) {real, imag} */,
  {32'hc54b4993, 32'h00000000} /* (25, 26, 0) {real, imag} */,
  {32'hc51a50b5, 32'h43d3fe31} /* (25, 25, 31) {real, imag} */,
  {32'h443ca530, 32'h43023fdc} /* (25, 25, 30) {real, imag} */,
  {32'hc12db634, 32'h42d03591} /* (25, 25, 29) {real, imag} */,
  {32'hc33db77a, 32'hc27ddc5b} /* (25, 25, 28) {real, imag} */,
  {32'h43580b20, 32'h41d3ee94} /* (25, 25, 27) {real, imag} */,
  {32'hbff68220, 32'hc13fe390} /* (25, 25, 26) {real, imag} */,
  {32'hc26b6e22, 32'h41c40c88} /* (25, 25, 25) {real, imag} */,
  {32'h424b405f, 32'h4227a7d0} /* (25, 25, 24) {real, imag} */,
  {32'h412aede6, 32'hc29eb650} /* (25, 25, 23) {real, imag} */,
  {32'h414ebed0, 32'h40dd6736} /* (25, 25, 22) {real, imag} */,
  {32'hc110d0a0, 32'hc2312db0} /* (25, 25, 21) {real, imag} */,
  {32'hc2bc66b2, 32'hc2964198} /* (25, 25, 20) {real, imag} */,
  {32'hc21f2b3e, 32'h429fe008} /* (25, 25, 19) {real, imag} */,
  {32'h42eec893, 32'hc242ac86} /* (25, 25, 18) {real, imag} */,
  {32'hc25f3fb1, 32'h426ce338} /* (25, 25, 17) {real, imag} */,
  {32'h423227d3, 32'h00000000} /* (25, 25, 16) {real, imag} */,
  {32'hc25f3fb1, 32'hc26ce338} /* (25, 25, 15) {real, imag} */,
  {32'h42eec893, 32'h4242ac86} /* (25, 25, 14) {real, imag} */,
  {32'hc21f2b3e, 32'hc29fe008} /* (25, 25, 13) {real, imag} */,
  {32'hc2bc66b2, 32'h42964198} /* (25, 25, 12) {real, imag} */,
  {32'hc110d0a0, 32'h42312db0} /* (25, 25, 11) {real, imag} */,
  {32'h414ebed0, 32'hc0dd6736} /* (25, 25, 10) {real, imag} */,
  {32'h412aede6, 32'h429eb650} /* (25, 25, 9) {real, imag} */,
  {32'h424b405f, 32'hc227a7d0} /* (25, 25, 8) {real, imag} */,
  {32'hc26b6e22, 32'hc1c40c88} /* (25, 25, 7) {real, imag} */,
  {32'hbff68220, 32'h413fe390} /* (25, 25, 6) {real, imag} */,
  {32'h43580b20, 32'hc1d3ee94} /* (25, 25, 5) {real, imag} */,
  {32'hc33db77a, 32'h427ddc5b} /* (25, 25, 4) {real, imag} */,
  {32'hc12db634, 32'hc2d03591} /* (25, 25, 3) {real, imag} */,
  {32'h443ca530, 32'hc3023fdc} /* (25, 25, 2) {real, imag} */,
  {32'hc51a50b5, 32'hc3d3fe31} /* (25, 25, 1) {real, imag} */,
  {32'hc5391734, 32'h00000000} /* (25, 25, 0) {real, imag} */,
  {32'hc50a7fde, 32'h43a08ec8} /* (25, 24, 31) {real, imag} */,
  {32'h4432013a, 32'hc1075d10} /* (25, 24, 30) {real, imag} */,
  {32'hc2d4405c, 32'hc03ccdb0} /* (25, 24, 29) {real, imag} */,
  {32'hc3362e9b, 32'hc2dd0065} /* (25, 24, 28) {real, imag} */,
  {32'h4345d0cd, 32'h4248c136} /* (25, 24, 27) {real, imag} */,
  {32'hc2730c21, 32'h40c8f920} /* (25, 24, 26) {real, imag} */,
  {32'h427fced0, 32'h3f61cc80} /* (25, 24, 25) {real, imag} */,
  {32'h41a34327, 32'hc2961af0} /* (25, 24, 24) {real, imag} */,
  {32'h40a7fe38, 32'hc1249ed2} /* (25, 24, 23) {real, imag} */,
  {32'hc278bbdb, 32'h42035de8} /* (25, 24, 22) {real, imag} */,
  {32'h4260fe0e, 32'hc2654026} /* (25, 24, 21) {real, imag} */,
  {32'h419bbe7b, 32'hc2d24d4e} /* (25, 24, 20) {real, imag} */,
  {32'h407f7320, 32'hc154d06a} /* (25, 24, 19) {real, imag} */,
  {32'h41ef9abc, 32'h416f54ac} /* (25, 24, 18) {real, imag} */,
  {32'h40878b20, 32'hc129b822} /* (25, 24, 17) {real, imag} */,
  {32'h42070e08, 32'h00000000} /* (25, 24, 16) {real, imag} */,
  {32'h40878b20, 32'h4129b822} /* (25, 24, 15) {real, imag} */,
  {32'h41ef9abc, 32'hc16f54ac} /* (25, 24, 14) {real, imag} */,
  {32'h407f7320, 32'h4154d06a} /* (25, 24, 13) {real, imag} */,
  {32'h419bbe7b, 32'h42d24d4e} /* (25, 24, 12) {real, imag} */,
  {32'h4260fe0e, 32'h42654026} /* (25, 24, 11) {real, imag} */,
  {32'hc278bbdb, 32'hc2035de8} /* (25, 24, 10) {real, imag} */,
  {32'h40a7fe38, 32'h41249ed2} /* (25, 24, 9) {real, imag} */,
  {32'h41a34327, 32'h42961af0} /* (25, 24, 8) {real, imag} */,
  {32'h427fced0, 32'hbf61cc80} /* (25, 24, 7) {real, imag} */,
  {32'hc2730c21, 32'hc0c8f920} /* (25, 24, 6) {real, imag} */,
  {32'h4345d0cd, 32'hc248c136} /* (25, 24, 5) {real, imag} */,
  {32'hc3362e9b, 32'h42dd0065} /* (25, 24, 4) {real, imag} */,
  {32'hc2d4405c, 32'h403ccdb0} /* (25, 24, 3) {real, imag} */,
  {32'h4432013a, 32'h41075d10} /* (25, 24, 2) {real, imag} */,
  {32'hc50a7fde, 32'hc3a08ec8} /* (25, 24, 1) {real, imag} */,
  {32'hc525242a, 32'h00000000} /* (25, 24, 0) {real, imag} */,
  {32'hc500cca2, 32'h439dabba} /* (25, 23, 31) {real, imag} */,
  {32'h443d60f9, 32'hc22dc232} /* (25, 23, 30) {real, imag} */,
  {32'hc22b8b86, 32'hc2bdfe11} /* (25, 23, 29) {real, imag} */,
  {32'hc1a1437a, 32'hc1eb9969} /* (25, 23, 28) {real, imag} */,
  {32'h4303177b, 32'h42ac4fea} /* (25, 23, 27) {real, imag} */,
  {32'hc2c416ff, 32'hc2e9aa46} /* (25, 23, 26) {real, imag} */,
  {32'hc2e84aae, 32'hc2145216} /* (25, 23, 25) {real, imag} */,
  {32'h4282fc14, 32'hc3247295} /* (25, 23, 24) {real, imag} */,
  {32'h3fb51ad0, 32'hc309b8b6} /* (25, 23, 23) {real, imag} */,
  {32'hc31c78ac, 32'h4245f62e} /* (25, 23, 22) {real, imag} */,
  {32'h42d1222c, 32'hc03b2ac0} /* (25, 23, 21) {real, imag} */,
  {32'hc18938b2, 32'hc11e89e5} /* (25, 23, 20) {real, imag} */,
  {32'h41fe8f4b, 32'hc2526232} /* (25, 23, 19) {real, imag} */,
  {32'hc1d6adf7, 32'h42969464} /* (25, 23, 18) {real, imag} */,
  {32'h42123fa2, 32'h4285d482} /* (25, 23, 17) {real, imag} */,
  {32'h419eb672, 32'h00000000} /* (25, 23, 16) {real, imag} */,
  {32'h42123fa2, 32'hc285d482} /* (25, 23, 15) {real, imag} */,
  {32'hc1d6adf7, 32'hc2969464} /* (25, 23, 14) {real, imag} */,
  {32'h41fe8f4b, 32'h42526232} /* (25, 23, 13) {real, imag} */,
  {32'hc18938b2, 32'h411e89e5} /* (25, 23, 12) {real, imag} */,
  {32'h42d1222c, 32'h403b2ac0} /* (25, 23, 11) {real, imag} */,
  {32'hc31c78ac, 32'hc245f62e} /* (25, 23, 10) {real, imag} */,
  {32'h3fb51ad0, 32'h4309b8b6} /* (25, 23, 9) {real, imag} */,
  {32'h4282fc14, 32'h43247295} /* (25, 23, 8) {real, imag} */,
  {32'hc2e84aae, 32'h42145216} /* (25, 23, 7) {real, imag} */,
  {32'hc2c416ff, 32'h42e9aa46} /* (25, 23, 6) {real, imag} */,
  {32'h4303177b, 32'hc2ac4fea} /* (25, 23, 5) {real, imag} */,
  {32'hc1a1437a, 32'h41eb9969} /* (25, 23, 4) {real, imag} */,
  {32'hc22b8b86, 32'h42bdfe11} /* (25, 23, 3) {real, imag} */,
  {32'h443d60f9, 32'h422dc232} /* (25, 23, 2) {real, imag} */,
  {32'hc500cca2, 32'hc39dabba} /* (25, 23, 1) {real, imag} */,
  {32'hc5073a84, 32'h00000000} /* (25, 23, 0) {real, imag} */,
  {32'hc4d3ca33, 32'h4338b5ad} /* (25, 22, 31) {real, imag} */,
  {32'h44290569, 32'hc2ef4ad7} /* (25, 22, 30) {real, imag} */,
  {32'h42894273, 32'h423b1076} /* (25, 22, 29) {real, imag} */,
  {32'hc2eff18f, 32'h42f7fa28} /* (25, 22, 28) {real, imag} */,
  {32'h433ad70a, 32'hc005f370} /* (25, 22, 27) {real, imag} */,
  {32'hc2090a14, 32'h42676af6} /* (25, 22, 26) {real, imag} */,
  {32'hc15eb0a2, 32'hc113b21c} /* (25, 22, 25) {real, imag} */,
  {32'h40a1498a, 32'hc129e730} /* (25, 22, 24) {real, imag} */,
  {32'h41af8ab9, 32'h42474d02} /* (25, 22, 23) {real, imag} */,
  {32'hc1058d50, 32'h4207ecc4} /* (25, 22, 22) {real, imag} */,
  {32'h40fc6458, 32'h42831f5e} /* (25, 22, 21) {real, imag} */,
  {32'hc01d97bc, 32'hc121181f} /* (25, 22, 20) {real, imag} */,
  {32'hc1d76e2c, 32'h42a2ada4} /* (25, 22, 19) {real, imag} */,
  {32'hc0c57a9b, 32'hc323da24} /* (25, 22, 18) {real, imag} */,
  {32'hbf97ad80, 32'hc211b12f} /* (25, 22, 17) {real, imag} */,
  {32'hc1baf0e2, 32'h00000000} /* (25, 22, 16) {real, imag} */,
  {32'hbf97ad80, 32'h4211b12f} /* (25, 22, 15) {real, imag} */,
  {32'hc0c57a9b, 32'h4323da24} /* (25, 22, 14) {real, imag} */,
  {32'hc1d76e2c, 32'hc2a2ada4} /* (25, 22, 13) {real, imag} */,
  {32'hc01d97bc, 32'h4121181f} /* (25, 22, 12) {real, imag} */,
  {32'h40fc6458, 32'hc2831f5e} /* (25, 22, 11) {real, imag} */,
  {32'hc1058d50, 32'hc207ecc4} /* (25, 22, 10) {real, imag} */,
  {32'h41af8ab9, 32'hc2474d02} /* (25, 22, 9) {real, imag} */,
  {32'h40a1498a, 32'h4129e730} /* (25, 22, 8) {real, imag} */,
  {32'hc15eb0a2, 32'h4113b21c} /* (25, 22, 7) {real, imag} */,
  {32'hc2090a14, 32'hc2676af6} /* (25, 22, 6) {real, imag} */,
  {32'h433ad70a, 32'h4005f370} /* (25, 22, 5) {real, imag} */,
  {32'hc2eff18f, 32'hc2f7fa28} /* (25, 22, 4) {real, imag} */,
  {32'h42894273, 32'hc23b1076} /* (25, 22, 3) {real, imag} */,
  {32'h44290569, 32'h42ef4ad7} /* (25, 22, 2) {real, imag} */,
  {32'hc4d3ca33, 32'hc338b5ad} /* (25, 22, 1) {real, imag} */,
  {32'hc4c08995, 32'h00000000} /* (25, 22, 0) {real, imag} */,
  {32'hc4557486, 32'h4225b850} /* (25, 21, 31) {real, imag} */,
  {32'h43e0308b, 32'h41f0a5d8} /* (25, 21, 30) {real, imag} */,
  {32'h419d84d8, 32'h4388aec2} /* (25, 21, 29) {real, imag} */,
  {32'hc33a9a70, 32'hc2b1bfa8} /* (25, 21, 28) {real, imag} */,
  {32'h42d72307, 32'hc27d84cc} /* (25, 21, 27) {real, imag} */,
  {32'h42ab7502, 32'h431f42fd} /* (25, 21, 26) {real, imag} */,
  {32'hc2ae99bc, 32'h4196d5ae} /* (25, 21, 25) {real, imag} */,
  {32'h41ff9706, 32'h41feaae8} /* (25, 21, 24) {real, imag} */,
  {32'h42f4255e, 32'hc1251810} /* (25, 21, 23) {real, imag} */,
  {32'h3fdbcf10, 32'hc00774bc} /* (25, 21, 22) {real, imag} */,
  {32'h42ae404c, 32'hc2dd4d40} /* (25, 21, 21) {real, imag} */,
  {32'h414506f4, 32'hc0ec3b1c} /* (25, 21, 20) {real, imag} */,
  {32'h4253047e, 32'hc14ebf40} /* (25, 21, 19) {real, imag} */,
  {32'hc2c838d1, 32'hbfa2d210} /* (25, 21, 18) {real, imag} */,
  {32'h426fe918, 32'hc24e005a} /* (25, 21, 17) {real, imag} */,
  {32'h430e407e, 32'h00000000} /* (25, 21, 16) {real, imag} */,
  {32'h426fe918, 32'h424e005a} /* (25, 21, 15) {real, imag} */,
  {32'hc2c838d1, 32'h3fa2d210} /* (25, 21, 14) {real, imag} */,
  {32'h4253047e, 32'h414ebf40} /* (25, 21, 13) {real, imag} */,
  {32'h414506f4, 32'h40ec3b1c} /* (25, 21, 12) {real, imag} */,
  {32'h42ae404c, 32'h42dd4d40} /* (25, 21, 11) {real, imag} */,
  {32'h3fdbcf10, 32'h400774bc} /* (25, 21, 10) {real, imag} */,
  {32'h42f4255e, 32'h41251810} /* (25, 21, 9) {real, imag} */,
  {32'h41ff9706, 32'hc1feaae8} /* (25, 21, 8) {real, imag} */,
  {32'hc2ae99bc, 32'hc196d5ae} /* (25, 21, 7) {real, imag} */,
  {32'h42ab7502, 32'hc31f42fd} /* (25, 21, 6) {real, imag} */,
  {32'h42d72307, 32'h427d84cc} /* (25, 21, 5) {real, imag} */,
  {32'hc33a9a70, 32'h42b1bfa8} /* (25, 21, 4) {real, imag} */,
  {32'h419d84d8, 32'hc388aec2} /* (25, 21, 3) {real, imag} */,
  {32'h43e0308b, 32'hc1f0a5d8} /* (25, 21, 2) {real, imag} */,
  {32'hc4557486, 32'hc225b850} /* (25, 21, 1) {real, imag} */,
  {32'hc44d75e1, 32'h00000000} /* (25, 21, 0) {real, imag} */,
  {32'h43a540c3, 32'hc2f9a600} /* (25, 20, 31) {real, imag} */,
  {32'hc3572a02, 32'h42de6b47} /* (25, 20, 30) {real, imag} */,
  {32'h42937ad7, 32'h4221f3f1} /* (25, 20, 29) {real, imag} */,
  {32'h40f7b6d0, 32'hc3246f21} /* (25, 20, 28) {real, imag} */,
  {32'hbedf2880, 32'h4297f18c} /* (25, 20, 27) {real, imag} */,
  {32'h42dc5198, 32'h435421e4} /* (25, 20, 26) {real, imag} */,
  {32'h423ae675, 32'hc28815ac} /* (25, 20, 25) {real, imag} */,
  {32'hc15c7088, 32'h428cc6e6} /* (25, 20, 24) {real, imag} */,
  {32'h40b1ca58, 32'hc25eeb8a} /* (25, 20, 23) {real, imag} */,
  {32'h428b096c, 32'h4270818c} /* (25, 20, 22) {real, imag} */,
  {32'h4268395e, 32'h423eb97a} /* (25, 20, 21) {real, imag} */,
  {32'h410de50c, 32'h41d1267c} /* (25, 20, 20) {real, imag} */,
  {32'hc1d547e7, 32'h42081c3a} /* (25, 20, 19) {real, imag} */,
  {32'hc264c3cf, 32'h40f25608} /* (25, 20, 18) {real, imag} */,
  {32'hc1aa032c, 32'hc2d62c29} /* (25, 20, 17) {real, imag} */,
  {32'h419e476e, 32'h00000000} /* (25, 20, 16) {real, imag} */,
  {32'hc1aa032c, 32'h42d62c29} /* (25, 20, 15) {real, imag} */,
  {32'hc264c3cf, 32'hc0f25608} /* (25, 20, 14) {real, imag} */,
  {32'hc1d547e7, 32'hc2081c3a} /* (25, 20, 13) {real, imag} */,
  {32'h410de50c, 32'hc1d1267c} /* (25, 20, 12) {real, imag} */,
  {32'h4268395e, 32'hc23eb97a} /* (25, 20, 11) {real, imag} */,
  {32'h428b096c, 32'hc270818c} /* (25, 20, 10) {real, imag} */,
  {32'h40b1ca58, 32'h425eeb8a} /* (25, 20, 9) {real, imag} */,
  {32'hc15c7088, 32'hc28cc6e6} /* (25, 20, 8) {real, imag} */,
  {32'h423ae675, 32'h428815ac} /* (25, 20, 7) {real, imag} */,
  {32'h42dc5198, 32'hc35421e4} /* (25, 20, 6) {real, imag} */,
  {32'hbedf2880, 32'hc297f18c} /* (25, 20, 5) {real, imag} */,
  {32'h40f7b6d0, 32'h43246f21} /* (25, 20, 4) {real, imag} */,
  {32'h42937ad7, 32'hc221f3f1} /* (25, 20, 3) {real, imag} */,
  {32'hc3572a02, 32'hc2de6b47} /* (25, 20, 2) {real, imag} */,
  {32'h43a540c3, 32'h42f9a600} /* (25, 20, 1) {real, imag} */,
  {32'h436e773c, 32'h00000000} /* (25, 20, 0) {real, imag} */,
  {32'h44501dd3, 32'hc328dd9a} /* (25, 19, 31) {real, imag} */,
  {32'hc3dbadfc, 32'hc214cfd2} /* (25, 19, 30) {real, imag} */,
  {32'h41808e78, 32'hc2a149fa} /* (25, 19, 29) {real, imag} */,
  {32'h43176daf, 32'hc2dda6a6} /* (25, 19, 28) {real, imag} */,
  {32'hc2e7492a, 32'h430e09be} /* (25, 19, 27) {real, imag} */,
  {32'h428a17b4, 32'hc16b9adc} /* (25, 19, 26) {real, imag} */,
  {32'h42cc416a, 32'hc27984d7} /* (25, 19, 25) {real, imag} */,
  {32'hc2f68fe1, 32'hc1c23691} /* (25, 19, 24) {real, imag} */,
  {32'h42033af6, 32'h3f85dbe0} /* (25, 19, 23) {real, imag} */,
  {32'h42a99394, 32'h4215d99c} /* (25, 19, 22) {real, imag} */,
  {32'hc2b23ee4, 32'h42a34434} /* (25, 19, 21) {real, imag} */,
  {32'hc12d9556, 32'hc1ffeea3} /* (25, 19, 20) {real, imag} */,
  {32'h41edb574, 32'hc1d1cf24} /* (25, 19, 19) {real, imag} */,
  {32'hc152a79e, 32'hc00ea40c} /* (25, 19, 18) {real, imag} */,
  {32'h413a6cb2, 32'hc136e4a6} /* (25, 19, 17) {real, imag} */,
  {32'hc29f6069, 32'h00000000} /* (25, 19, 16) {real, imag} */,
  {32'h413a6cb2, 32'h4136e4a6} /* (25, 19, 15) {real, imag} */,
  {32'hc152a79e, 32'h400ea40c} /* (25, 19, 14) {real, imag} */,
  {32'h41edb574, 32'h41d1cf24} /* (25, 19, 13) {real, imag} */,
  {32'hc12d9556, 32'h41ffeea3} /* (25, 19, 12) {real, imag} */,
  {32'hc2b23ee4, 32'hc2a34434} /* (25, 19, 11) {real, imag} */,
  {32'h42a99394, 32'hc215d99c} /* (25, 19, 10) {real, imag} */,
  {32'h42033af6, 32'hbf85dbe0} /* (25, 19, 9) {real, imag} */,
  {32'hc2f68fe1, 32'h41c23691} /* (25, 19, 8) {real, imag} */,
  {32'h42cc416a, 32'h427984d7} /* (25, 19, 7) {real, imag} */,
  {32'h428a17b4, 32'h416b9adc} /* (25, 19, 6) {real, imag} */,
  {32'hc2e7492a, 32'hc30e09be} /* (25, 19, 5) {real, imag} */,
  {32'h43176daf, 32'h42dda6a6} /* (25, 19, 4) {real, imag} */,
  {32'h41808e78, 32'h42a149fa} /* (25, 19, 3) {real, imag} */,
  {32'hc3dbadfc, 32'h4214cfd2} /* (25, 19, 2) {real, imag} */,
  {32'h44501dd3, 32'h4328dd9a} /* (25, 19, 1) {real, imag} */,
  {32'h4440d512, 32'h00000000} /* (25, 19, 0) {real, imag} */,
  {32'h44a10cca, 32'hc2ca50c8} /* (25, 18, 31) {real, imag} */,
  {32'hc407810a, 32'h420136aa} /* (25, 18, 30) {real, imag} */,
  {32'hc0192d50, 32'hc0e3e038} /* (25, 18, 29) {real, imag} */,
  {32'h435d357e, 32'hc28fba7c} /* (25, 18, 28) {real, imag} */,
  {32'h4103169c, 32'h42a4c8e5} /* (25, 18, 27) {real, imag} */,
  {32'h41655bee, 32'h4051da28} /* (25, 18, 26) {real, imag} */,
  {32'hc1b7773e, 32'hc093f218} /* (25, 18, 25) {real, imag} */,
  {32'hc2980f82, 32'hc28443d4} /* (25, 18, 24) {real, imag} */,
  {32'hc3118a32, 32'hc1659938} /* (25, 18, 23) {real, imag} */,
  {32'hc2adedf4, 32'hc2193cf0} /* (25, 18, 22) {real, imag} */,
  {32'hc2296d15, 32'hc113498c} /* (25, 18, 21) {real, imag} */,
  {32'h40d8171c, 32'h42155d6a} /* (25, 18, 20) {real, imag} */,
  {32'hc23bfe29, 32'hc2a8b482} /* (25, 18, 19) {real, imag} */,
  {32'h4226b13b, 32'hc28394ec} /* (25, 18, 18) {real, imag} */,
  {32'h4124207e, 32'h4106daca} /* (25, 18, 17) {real, imag} */,
  {32'h4244df2f, 32'h00000000} /* (25, 18, 16) {real, imag} */,
  {32'h4124207e, 32'hc106daca} /* (25, 18, 15) {real, imag} */,
  {32'h4226b13b, 32'h428394ec} /* (25, 18, 14) {real, imag} */,
  {32'hc23bfe29, 32'h42a8b482} /* (25, 18, 13) {real, imag} */,
  {32'h40d8171c, 32'hc2155d6a} /* (25, 18, 12) {real, imag} */,
  {32'hc2296d15, 32'h4113498c} /* (25, 18, 11) {real, imag} */,
  {32'hc2adedf4, 32'h42193cf0} /* (25, 18, 10) {real, imag} */,
  {32'hc3118a32, 32'h41659938} /* (25, 18, 9) {real, imag} */,
  {32'hc2980f82, 32'h428443d4} /* (25, 18, 8) {real, imag} */,
  {32'hc1b7773e, 32'h4093f218} /* (25, 18, 7) {real, imag} */,
  {32'h41655bee, 32'hc051da28} /* (25, 18, 6) {real, imag} */,
  {32'h4103169c, 32'hc2a4c8e5} /* (25, 18, 5) {real, imag} */,
  {32'h435d357e, 32'h428fba7c} /* (25, 18, 4) {real, imag} */,
  {32'hc0192d50, 32'h40e3e038} /* (25, 18, 3) {real, imag} */,
  {32'hc407810a, 32'hc20136aa} /* (25, 18, 2) {real, imag} */,
  {32'h44a10cca, 32'h42ca50c8} /* (25, 18, 1) {real, imag} */,
  {32'h447a8d04, 32'h00000000} /* (25, 18, 0) {real, imag} */,
  {32'h44c39ba2, 32'hc34336e5} /* (25, 17, 31) {real, imag} */,
  {32'hc445f14a, 32'h42a120c6} /* (25, 17, 30) {real, imag} */,
  {32'hc29b7d5e, 32'hc26d0752} /* (25, 17, 29) {real, imag} */,
  {32'h435e4f30, 32'hc28d58f6} /* (25, 17, 28) {real, imag} */,
  {32'hc27b919d, 32'h42a43691} /* (25, 17, 27) {real, imag} */,
  {32'hc2011020, 32'h429dcb9a} /* (25, 17, 26) {real, imag} */,
  {32'hc2066fa4, 32'h412c1bfa} /* (25, 17, 25) {real, imag} */,
  {32'hc0e8be68, 32'hc29646ad} /* (25, 17, 24) {real, imag} */,
  {32'h407fdaf8, 32'hc1e5d194} /* (25, 17, 23) {real, imag} */,
  {32'hc13ee21f, 32'hc20afbfc} /* (25, 17, 22) {real, imag} */,
  {32'hc107efb0, 32'h426af270} /* (25, 17, 21) {real, imag} */,
  {32'h42306848, 32'hc27499b7} /* (25, 17, 20) {real, imag} */,
  {32'h4274a3dc, 32'hc245f596} /* (25, 17, 19) {real, imag} */,
  {32'h418029c8, 32'h41c915d7} /* (25, 17, 18) {real, imag} */,
  {32'hc17ffa56, 32'hc11a131c} /* (25, 17, 17) {real, imag} */,
  {32'hc1d47347, 32'h00000000} /* (25, 17, 16) {real, imag} */,
  {32'hc17ffa56, 32'h411a131c} /* (25, 17, 15) {real, imag} */,
  {32'h418029c8, 32'hc1c915d7} /* (25, 17, 14) {real, imag} */,
  {32'h4274a3dc, 32'h4245f596} /* (25, 17, 13) {real, imag} */,
  {32'h42306848, 32'h427499b7} /* (25, 17, 12) {real, imag} */,
  {32'hc107efb0, 32'hc26af270} /* (25, 17, 11) {real, imag} */,
  {32'hc13ee21f, 32'h420afbfc} /* (25, 17, 10) {real, imag} */,
  {32'h407fdaf8, 32'h41e5d194} /* (25, 17, 9) {real, imag} */,
  {32'hc0e8be68, 32'h429646ad} /* (25, 17, 8) {real, imag} */,
  {32'hc2066fa4, 32'hc12c1bfa} /* (25, 17, 7) {real, imag} */,
  {32'hc2011020, 32'hc29dcb9a} /* (25, 17, 6) {real, imag} */,
  {32'hc27b919d, 32'hc2a43691} /* (25, 17, 5) {real, imag} */,
  {32'h435e4f30, 32'h428d58f6} /* (25, 17, 4) {real, imag} */,
  {32'hc29b7d5e, 32'h426d0752} /* (25, 17, 3) {real, imag} */,
  {32'hc445f14a, 32'hc2a120c6} /* (25, 17, 2) {real, imag} */,
  {32'h44c39ba2, 32'h434336e5} /* (25, 17, 1) {real, imag} */,
  {32'h44a2e52d, 32'h00000000} /* (25, 17, 0) {real, imag} */,
  {32'h44ed3f81, 32'hc22ebb10} /* (25, 16, 31) {real, imag} */,
  {32'hc42810da, 32'h439bb818} /* (25, 16, 30) {real, imag} */,
  {32'hc3369933, 32'hc29bdc8c} /* (25, 16, 29) {real, imag} */,
  {32'h432dbb53, 32'hc32d734a} /* (25, 16, 28) {real, imag} */,
  {32'hc21fc86a, 32'h41e48eff} /* (25, 16, 27) {real, imag} */,
  {32'hc16c1af4, 32'h428fdf38} /* (25, 16, 26) {real, imag} */,
  {32'hc194a3cc, 32'h42b2415e} /* (25, 16, 25) {real, imag} */,
  {32'hc2cace42, 32'hc1d5061e} /* (25, 16, 24) {real, imag} */,
  {32'h42bf5dae, 32'hc2d6dcba} /* (25, 16, 23) {real, imag} */,
  {32'h430afe26, 32'hc29377c8} /* (25, 16, 22) {real, imag} */,
  {32'h41e3feb0, 32'h4154bbf4} /* (25, 16, 21) {real, imag} */,
  {32'hc2ba3fe3, 32'h425dea0a} /* (25, 16, 20) {real, imag} */,
  {32'hc116d99c, 32'h42e401ab} /* (25, 16, 19) {real, imag} */,
  {32'hc220b36c, 32'hc1556146} /* (25, 16, 18) {real, imag} */,
  {32'h42a988d6, 32'hc294e10c} /* (25, 16, 17) {real, imag} */,
  {32'h42a3991d, 32'h00000000} /* (25, 16, 16) {real, imag} */,
  {32'h42a988d6, 32'h4294e10c} /* (25, 16, 15) {real, imag} */,
  {32'hc220b36c, 32'h41556146} /* (25, 16, 14) {real, imag} */,
  {32'hc116d99c, 32'hc2e401ab} /* (25, 16, 13) {real, imag} */,
  {32'hc2ba3fe3, 32'hc25dea0a} /* (25, 16, 12) {real, imag} */,
  {32'h41e3feb0, 32'hc154bbf4} /* (25, 16, 11) {real, imag} */,
  {32'h430afe26, 32'h429377c8} /* (25, 16, 10) {real, imag} */,
  {32'h42bf5dae, 32'h42d6dcba} /* (25, 16, 9) {real, imag} */,
  {32'hc2cace42, 32'h41d5061e} /* (25, 16, 8) {real, imag} */,
  {32'hc194a3cc, 32'hc2b2415e} /* (25, 16, 7) {real, imag} */,
  {32'hc16c1af4, 32'hc28fdf38} /* (25, 16, 6) {real, imag} */,
  {32'hc21fc86a, 32'hc1e48eff} /* (25, 16, 5) {real, imag} */,
  {32'h432dbb53, 32'h432d734a} /* (25, 16, 4) {real, imag} */,
  {32'hc3369933, 32'h429bdc8c} /* (25, 16, 3) {real, imag} */,
  {32'hc42810da, 32'hc39bb818} /* (25, 16, 2) {real, imag} */,
  {32'h44ed3f81, 32'h422ebb10} /* (25, 16, 1) {real, imag} */,
  {32'h44aed6c8, 32'h00000000} /* (25, 16, 0) {real, imag} */,
  {32'h44e669fa, 32'hc1b0c298} /* (25, 15, 31) {real, imag} */,
  {32'hc4242b78, 32'h43281d5d} /* (25, 15, 30) {real, imag} */,
  {32'h42094f28, 32'hc21b8226} /* (25, 15, 29) {real, imag} */,
  {32'h40eb36f0, 32'hc312aecd} /* (25, 15, 28) {real, imag} */,
  {32'hc32e0995, 32'hbf87d540} /* (25, 15, 27) {real, imag} */,
  {32'hc1ddc088, 32'h4207a248} /* (25, 15, 26) {real, imag} */,
  {32'h42c1bb5c, 32'hc219846c} /* (25, 15, 25) {real, imag} */,
  {32'h41780ba4, 32'hc0fd1db0} /* (25, 15, 24) {real, imag} */,
  {32'hbff2e650, 32'hc12ab628} /* (25, 15, 23) {real, imag} */,
  {32'h4175dbfd, 32'hc100eff3} /* (25, 15, 22) {real, imag} */,
  {32'hc107b02c, 32'h420c4cf8} /* (25, 15, 21) {real, imag} */,
  {32'hc24fec3c, 32'hc2545899} /* (25, 15, 20) {real, imag} */,
  {32'hc232588c, 32'h422afe4a} /* (25, 15, 19) {real, imag} */,
  {32'h41ff6388, 32'hc0ba92fc} /* (25, 15, 18) {real, imag} */,
  {32'h41ba6047, 32'h414ad582} /* (25, 15, 17) {real, imag} */,
  {32'h42055eea, 32'h00000000} /* (25, 15, 16) {real, imag} */,
  {32'h41ba6047, 32'hc14ad582} /* (25, 15, 15) {real, imag} */,
  {32'h41ff6388, 32'h40ba92fc} /* (25, 15, 14) {real, imag} */,
  {32'hc232588c, 32'hc22afe4a} /* (25, 15, 13) {real, imag} */,
  {32'hc24fec3c, 32'h42545899} /* (25, 15, 12) {real, imag} */,
  {32'hc107b02c, 32'hc20c4cf8} /* (25, 15, 11) {real, imag} */,
  {32'h4175dbfd, 32'h4100eff3} /* (25, 15, 10) {real, imag} */,
  {32'hbff2e650, 32'h412ab628} /* (25, 15, 9) {real, imag} */,
  {32'h41780ba4, 32'h40fd1db0} /* (25, 15, 8) {real, imag} */,
  {32'h42c1bb5c, 32'h4219846c} /* (25, 15, 7) {real, imag} */,
  {32'hc1ddc088, 32'hc207a248} /* (25, 15, 6) {real, imag} */,
  {32'hc32e0995, 32'h3f87d540} /* (25, 15, 5) {real, imag} */,
  {32'h40eb36f0, 32'h4312aecd} /* (25, 15, 4) {real, imag} */,
  {32'h42094f28, 32'h421b8226} /* (25, 15, 3) {real, imag} */,
  {32'hc4242b78, 32'hc3281d5d} /* (25, 15, 2) {real, imag} */,
  {32'h44e669fa, 32'h41b0c298} /* (25, 15, 1) {real, imag} */,
  {32'h4491929b, 32'h00000000} /* (25, 15, 0) {real, imag} */,
  {32'h44deda42, 32'hc101b1c0} /* (25, 14, 31) {real, imag} */,
  {32'hc436137e, 32'h43164948} /* (25, 14, 30) {real, imag} */,
  {32'hc1bdb2f6, 32'hc235a6d9} /* (25, 14, 29) {real, imag} */,
  {32'h420a3184, 32'hc2aaf5a8} /* (25, 14, 28) {real, imag} */,
  {32'hc2b2cfd2, 32'h428c36af} /* (25, 14, 27) {real, imag} */,
  {32'h415404f8, 32'hc1312806} /* (25, 14, 26) {real, imag} */,
  {32'h42281637, 32'hc14404a8} /* (25, 14, 25) {real, imag} */,
  {32'hc14d74c0, 32'h402e3440} /* (25, 14, 24) {real, imag} */,
  {32'hc0154c20, 32'h419b0778} /* (25, 14, 23) {real, imag} */,
  {32'hc27ce399, 32'h428f405c} /* (25, 14, 22) {real, imag} */,
  {32'h42389ac3, 32'h41d57782} /* (25, 14, 21) {real, imag} */,
  {32'hc2556476, 32'hc09f163c} /* (25, 14, 20) {real, imag} */,
  {32'h41d1c31a, 32'hc205ca54} /* (25, 14, 19) {real, imag} */,
  {32'hc19d3d74, 32'h41a91957} /* (25, 14, 18) {real, imag} */,
  {32'hc23ab926, 32'hc1be9ee3} /* (25, 14, 17) {real, imag} */,
  {32'hc29534a0, 32'h00000000} /* (25, 14, 16) {real, imag} */,
  {32'hc23ab926, 32'h41be9ee3} /* (25, 14, 15) {real, imag} */,
  {32'hc19d3d74, 32'hc1a91957} /* (25, 14, 14) {real, imag} */,
  {32'h41d1c31a, 32'h4205ca54} /* (25, 14, 13) {real, imag} */,
  {32'hc2556476, 32'h409f163c} /* (25, 14, 12) {real, imag} */,
  {32'h42389ac3, 32'hc1d57782} /* (25, 14, 11) {real, imag} */,
  {32'hc27ce399, 32'hc28f405c} /* (25, 14, 10) {real, imag} */,
  {32'hc0154c20, 32'hc19b0778} /* (25, 14, 9) {real, imag} */,
  {32'hc14d74c0, 32'hc02e3440} /* (25, 14, 8) {real, imag} */,
  {32'h42281637, 32'h414404a8} /* (25, 14, 7) {real, imag} */,
  {32'h415404f8, 32'h41312806} /* (25, 14, 6) {real, imag} */,
  {32'hc2b2cfd2, 32'hc28c36af} /* (25, 14, 5) {real, imag} */,
  {32'h420a3184, 32'h42aaf5a8} /* (25, 14, 4) {real, imag} */,
  {32'hc1bdb2f6, 32'h4235a6d9} /* (25, 14, 3) {real, imag} */,
  {32'hc436137e, 32'hc3164948} /* (25, 14, 2) {real, imag} */,
  {32'h44deda42, 32'h4101b1c0} /* (25, 14, 1) {real, imag} */,
  {32'h446e84a4, 32'h00000000} /* (25, 14, 0) {real, imag} */,
  {32'h44ccf586, 32'h421e9b28} /* (25, 13, 31) {real, imag} */,
  {32'hc44a8096, 32'h431f4b84} /* (25, 13, 30) {real, imag} */,
  {32'hc250b650, 32'hc1871f1e} /* (25, 13, 29) {real, imag} */,
  {32'hc1c13210, 32'hc2e45b80} /* (25, 13, 28) {real, imag} */,
  {32'hc2c5af9e, 32'hc1b40144} /* (25, 13, 27) {real, imag} */,
  {32'hc24888f8, 32'h4132cc18} /* (25, 13, 26) {real, imag} */,
  {32'h43372d59, 32'hc1158864} /* (25, 13, 25) {real, imag} */,
  {32'hc2b37f07, 32'h4022ae10} /* (25, 13, 24) {real, imag} */,
  {32'h42835ec8, 32'hc19e5c84} /* (25, 13, 23) {real, imag} */,
  {32'hc1ec4022, 32'h41175e3a} /* (25, 13, 22) {real, imag} */,
  {32'hc28d2db4, 32'h42a7ebe0} /* (25, 13, 21) {real, imag} */,
  {32'hc24002bc, 32'h413c255a} /* (25, 13, 20) {real, imag} */,
  {32'h42828db8, 32'h41b5c198} /* (25, 13, 19) {real, imag} */,
  {32'h41770f60, 32'h3fc814f8} /* (25, 13, 18) {real, imag} */,
  {32'h423cb420, 32'hc1963679} /* (25, 13, 17) {real, imag} */,
  {32'h416d9748, 32'h00000000} /* (25, 13, 16) {real, imag} */,
  {32'h423cb420, 32'h41963679} /* (25, 13, 15) {real, imag} */,
  {32'h41770f60, 32'hbfc814f8} /* (25, 13, 14) {real, imag} */,
  {32'h42828db8, 32'hc1b5c198} /* (25, 13, 13) {real, imag} */,
  {32'hc24002bc, 32'hc13c255a} /* (25, 13, 12) {real, imag} */,
  {32'hc28d2db4, 32'hc2a7ebe0} /* (25, 13, 11) {real, imag} */,
  {32'hc1ec4022, 32'hc1175e3a} /* (25, 13, 10) {real, imag} */,
  {32'h42835ec8, 32'h419e5c84} /* (25, 13, 9) {real, imag} */,
  {32'hc2b37f07, 32'hc022ae10} /* (25, 13, 8) {real, imag} */,
  {32'h43372d59, 32'h41158864} /* (25, 13, 7) {real, imag} */,
  {32'hc24888f8, 32'hc132cc18} /* (25, 13, 6) {real, imag} */,
  {32'hc2c5af9e, 32'h41b40144} /* (25, 13, 5) {real, imag} */,
  {32'hc1c13210, 32'h42e45b80} /* (25, 13, 4) {real, imag} */,
  {32'hc250b650, 32'h41871f1e} /* (25, 13, 3) {real, imag} */,
  {32'hc44a8096, 32'hc31f4b84} /* (25, 13, 2) {real, imag} */,
  {32'h44ccf586, 32'hc21e9b28} /* (25, 13, 1) {real, imag} */,
  {32'h4489f4cb, 32'h00000000} /* (25, 13, 0) {real, imag} */,
  {32'h44a7e78d, 32'h43436ab0} /* (25, 12, 31) {real, imag} */,
  {32'hc43b368e, 32'hc11fb568} /* (25, 12, 30) {real, imag} */,
  {32'h412f3f78, 32'h40ef3b10} /* (25, 12, 29) {real, imag} */,
  {32'h431c49e6, 32'hc328c93d} /* (25, 12, 28) {real, imag} */,
  {32'hc2fa694a, 32'h417c1c70} /* (25, 12, 27) {real, imag} */,
  {32'hbe8c2980, 32'hc1ab359c} /* (25, 12, 26) {real, imag} */,
  {32'h42185d2b, 32'h41eb191a} /* (25, 12, 25) {real, imag} */,
  {32'hc2e204b3, 32'h42ff09d0} /* (25, 12, 24) {real, imag} */,
  {32'hc28eb9ee, 32'hc31f81a4} /* (25, 12, 23) {real, imag} */,
  {32'hc1479d90, 32'hc0995a40} /* (25, 12, 22) {real, imag} */,
  {32'hc314f41c, 32'h42c19ec7} /* (25, 12, 21) {real, imag} */,
  {32'hc2680109, 32'hc1be5148} /* (25, 12, 20) {real, imag} */,
  {32'h42005e00, 32'h41bad49b} /* (25, 12, 19) {real, imag} */,
  {32'hc127ae64, 32'h4288c0be} /* (25, 12, 18) {real, imag} */,
  {32'h41b973c8, 32'hc279c54a} /* (25, 12, 17) {real, imag} */,
  {32'h415b8c04, 32'h00000000} /* (25, 12, 16) {real, imag} */,
  {32'h41b973c8, 32'h4279c54a} /* (25, 12, 15) {real, imag} */,
  {32'hc127ae64, 32'hc288c0be} /* (25, 12, 14) {real, imag} */,
  {32'h42005e00, 32'hc1bad49b} /* (25, 12, 13) {real, imag} */,
  {32'hc2680109, 32'h41be5148} /* (25, 12, 12) {real, imag} */,
  {32'hc314f41c, 32'hc2c19ec7} /* (25, 12, 11) {real, imag} */,
  {32'hc1479d90, 32'h40995a40} /* (25, 12, 10) {real, imag} */,
  {32'hc28eb9ee, 32'h431f81a4} /* (25, 12, 9) {real, imag} */,
  {32'hc2e204b3, 32'hc2ff09d0} /* (25, 12, 8) {real, imag} */,
  {32'h42185d2b, 32'hc1eb191a} /* (25, 12, 7) {real, imag} */,
  {32'hbe8c2980, 32'h41ab359c} /* (25, 12, 6) {real, imag} */,
  {32'hc2fa694a, 32'hc17c1c70} /* (25, 12, 5) {real, imag} */,
  {32'h431c49e6, 32'h4328c93d} /* (25, 12, 4) {real, imag} */,
  {32'h412f3f78, 32'hc0ef3b10} /* (25, 12, 3) {real, imag} */,
  {32'hc43b368e, 32'h411fb568} /* (25, 12, 2) {real, imag} */,
  {32'h44a7e78d, 32'hc3436ab0} /* (25, 12, 1) {real, imag} */,
  {32'h443eb545, 32'h00000000} /* (25, 12, 0) {real, imag} */,
  {32'h443c549e, 32'h439e96ea} /* (25, 11, 31) {real, imag} */,
  {32'hc410c71c, 32'h42223f60} /* (25, 11, 30) {real, imag} */,
  {32'hc11180fd, 32'h40983020} /* (25, 11, 29) {real, imag} */,
  {32'h438af096, 32'hc389c1f2} /* (25, 11, 28) {real, imag} */,
  {32'hc1f6d574, 32'h43339d82} /* (25, 11, 27) {real, imag} */,
  {32'hc209918d, 32'h41866608} /* (25, 11, 26) {real, imag} */,
  {32'hbe1f8100, 32'h422ac431} /* (25, 11, 25) {real, imag} */,
  {32'h4214c1b9, 32'hc0d379a0} /* (25, 11, 24) {real, imag} */,
  {32'hc1c421ae, 32'h422fd960} /* (25, 11, 23) {real, imag} */,
  {32'h427b6bfc, 32'hc10b2655} /* (25, 11, 22) {real, imag} */,
  {32'hc2e071c4, 32'h426be768} /* (25, 11, 21) {real, imag} */,
  {32'h41a94470, 32'h41e559df} /* (25, 11, 20) {real, imag} */,
  {32'hc00f15f8, 32'hc0f5c470} /* (25, 11, 19) {real, imag} */,
  {32'h41475a60, 32'h426036f2} /* (25, 11, 18) {real, imag} */,
  {32'hc17306d0, 32'h4193e3ab} /* (25, 11, 17) {real, imag} */,
  {32'h41d79996, 32'h00000000} /* (25, 11, 16) {real, imag} */,
  {32'hc17306d0, 32'hc193e3ab} /* (25, 11, 15) {real, imag} */,
  {32'h41475a60, 32'hc26036f2} /* (25, 11, 14) {real, imag} */,
  {32'hc00f15f8, 32'h40f5c470} /* (25, 11, 13) {real, imag} */,
  {32'h41a94470, 32'hc1e559df} /* (25, 11, 12) {real, imag} */,
  {32'hc2e071c4, 32'hc26be768} /* (25, 11, 11) {real, imag} */,
  {32'h427b6bfc, 32'h410b2655} /* (25, 11, 10) {real, imag} */,
  {32'hc1c421ae, 32'hc22fd960} /* (25, 11, 9) {real, imag} */,
  {32'h4214c1b9, 32'h40d379a0} /* (25, 11, 8) {real, imag} */,
  {32'hbe1f8100, 32'hc22ac431} /* (25, 11, 7) {real, imag} */,
  {32'hc209918d, 32'hc1866608} /* (25, 11, 6) {real, imag} */,
  {32'hc1f6d574, 32'hc3339d82} /* (25, 11, 5) {real, imag} */,
  {32'h438af096, 32'h4389c1f2} /* (25, 11, 4) {real, imag} */,
  {32'hc11180fd, 32'hc0983020} /* (25, 11, 3) {real, imag} */,
  {32'hc410c71c, 32'hc2223f60} /* (25, 11, 2) {real, imag} */,
  {32'h443c549e, 32'hc39e96ea} /* (25, 11, 1) {real, imag} */,
  {32'h43c542d2, 32'h00000000} /* (25, 11, 0) {real, imag} */,
  {32'hc4050f12, 32'h440d852c} /* (25, 10, 31) {real, imag} */,
  {32'hc21ac590, 32'h418b4054} /* (25, 10, 30) {real, imag} */,
  {32'hc2158c3e, 32'hc301748c} /* (25, 10, 29) {real, imag} */,
  {32'h42f7fc51, 32'hc291609c} /* (25, 10, 28) {real, imag} */,
  {32'hc17e5f60, 32'hc2d8d3f0} /* (25, 10, 27) {real, imag} */,
  {32'h4212ec60, 32'h41d21759} /* (25, 10, 26) {real, imag} */,
  {32'hc28aef2e, 32'h41610924} /* (25, 10, 25) {real, imag} */,
  {32'hc194d028, 32'hc33b3eae} /* (25, 10, 24) {real, imag} */,
  {32'h412d6b36, 32'hc2bffa63} /* (25, 10, 23) {real, imag} */,
  {32'hc2869e3f, 32'h426899d4} /* (25, 10, 22) {real, imag} */,
  {32'hc2972fca, 32'hc246f238} /* (25, 10, 21) {real, imag} */,
  {32'hc1bd8b9e, 32'hc15d378f} /* (25, 10, 20) {real, imag} */,
  {32'h423eb314, 32'hc2f1c8a8} /* (25, 10, 19) {real, imag} */,
  {32'h41a14ed0, 32'h41c23868} /* (25, 10, 18) {real, imag} */,
  {32'h42a0f19d, 32'h42c03a50} /* (25, 10, 17) {real, imag} */,
  {32'hc21bbc51, 32'h00000000} /* (25, 10, 16) {real, imag} */,
  {32'h42a0f19d, 32'hc2c03a50} /* (25, 10, 15) {real, imag} */,
  {32'h41a14ed0, 32'hc1c23868} /* (25, 10, 14) {real, imag} */,
  {32'h423eb314, 32'h42f1c8a8} /* (25, 10, 13) {real, imag} */,
  {32'hc1bd8b9e, 32'h415d378f} /* (25, 10, 12) {real, imag} */,
  {32'hc2972fca, 32'h4246f238} /* (25, 10, 11) {real, imag} */,
  {32'hc2869e3f, 32'hc26899d4} /* (25, 10, 10) {real, imag} */,
  {32'h412d6b36, 32'h42bffa63} /* (25, 10, 9) {real, imag} */,
  {32'hc194d028, 32'h433b3eae} /* (25, 10, 8) {real, imag} */,
  {32'hc28aef2e, 32'hc1610924} /* (25, 10, 7) {real, imag} */,
  {32'h4212ec60, 32'hc1d21759} /* (25, 10, 6) {real, imag} */,
  {32'hc17e5f60, 32'h42d8d3f0} /* (25, 10, 5) {real, imag} */,
  {32'h42f7fc51, 32'h4291609c} /* (25, 10, 4) {real, imag} */,
  {32'hc2158c3e, 32'h4301748c} /* (25, 10, 3) {real, imag} */,
  {32'hc21ac590, 32'hc18b4054} /* (25, 10, 2) {real, imag} */,
  {32'hc4050f12, 32'hc40d852c} /* (25, 10, 1) {real, imag} */,
  {32'hc414fe9e, 32'h00000000} /* (25, 10, 0) {real, imag} */,
  {32'hc498875b, 32'h442f5b2e} /* (25, 9, 31) {real, imag} */,
  {32'h4382e2e8, 32'hc2caa217} /* (25, 9, 30) {real, imag} */,
  {32'h424abd54, 32'hc242ebee} /* (25, 9, 29) {real, imag} */,
  {32'hc1af85f2, 32'hc27978bc} /* (25, 9, 28) {real, imag} */,
  {32'h427c523f, 32'hc2f47982} /* (25, 9, 27) {real, imag} */,
  {32'hc2634a7e, 32'h3ee90100} /* (25, 9, 26) {real, imag} */,
  {32'hc15361a0, 32'h42873554} /* (25, 9, 25) {real, imag} */,
  {32'hc1a67ca8, 32'hc282ac54} /* (25, 9, 24) {real, imag} */,
  {32'h42015b90, 32'hc257d678} /* (25, 9, 23) {real, imag} */,
  {32'h421b822a, 32'hbfd82a90} /* (25, 9, 22) {real, imag} */,
  {32'h4211a99f, 32'hc2a9d15b} /* (25, 9, 21) {real, imag} */,
  {32'hc2919826, 32'h4192eb2a} /* (25, 9, 20) {real, imag} */,
  {32'hc1774cea, 32'h3f2734e0} /* (25, 9, 19) {real, imag} */,
  {32'h425e0442, 32'hc1b8783f} /* (25, 9, 18) {real, imag} */,
  {32'hc19f7720, 32'hc0e5c684} /* (25, 9, 17) {real, imag} */,
  {32'h420bfa71, 32'h00000000} /* (25, 9, 16) {real, imag} */,
  {32'hc19f7720, 32'h40e5c684} /* (25, 9, 15) {real, imag} */,
  {32'h425e0442, 32'h41b8783f} /* (25, 9, 14) {real, imag} */,
  {32'hc1774cea, 32'hbf2734e0} /* (25, 9, 13) {real, imag} */,
  {32'hc2919826, 32'hc192eb2a} /* (25, 9, 12) {real, imag} */,
  {32'h4211a99f, 32'h42a9d15b} /* (25, 9, 11) {real, imag} */,
  {32'h421b822a, 32'h3fd82a90} /* (25, 9, 10) {real, imag} */,
  {32'h42015b90, 32'h4257d678} /* (25, 9, 9) {real, imag} */,
  {32'hc1a67ca8, 32'h4282ac54} /* (25, 9, 8) {real, imag} */,
  {32'hc15361a0, 32'hc2873554} /* (25, 9, 7) {real, imag} */,
  {32'hc2634a7e, 32'hbee90100} /* (25, 9, 6) {real, imag} */,
  {32'h427c523f, 32'h42f47982} /* (25, 9, 5) {real, imag} */,
  {32'hc1af85f2, 32'h427978bc} /* (25, 9, 4) {real, imag} */,
  {32'h424abd54, 32'h4242ebee} /* (25, 9, 3) {real, imag} */,
  {32'h4382e2e8, 32'h42caa217} /* (25, 9, 2) {real, imag} */,
  {32'hc498875b, 32'hc42f5b2e} /* (25, 9, 1) {real, imag} */,
  {32'hc4ae249c, 32'h00000000} /* (25, 9, 0) {real, imag} */,
  {32'hc4c5deb3, 32'h44569bae} /* (25, 8, 31) {real, imag} */,
  {32'h43cbae23, 32'hc30589df} /* (25, 8, 30) {real, imag} */,
  {32'h420200f7, 32'hc1abc3e6} /* (25, 8, 29) {real, imag} */,
  {32'hc2a8870e, 32'h4194deac} /* (25, 8, 28) {real, imag} */,
  {32'h4201ab4c, 32'hc25e7e7e} /* (25, 8, 27) {real, imag} */,
  {32'hc265d837, 32'hc2d7a465} /* (25, 8, 26) {real, imag} */,
  {32'hc15ee60e, 32'hc29d5b88} /* (25, 8, 25) {real, imag} */,
  {32'hc02618e8, 32'hc31cdbf0} /* (25, 8, 24) {real, imag} */,
  {32'hc2800664, 32'hc1bb48fb} /* (25, 8, 23) {real, imag} */,
  {32'hc2744fcf, 32'h4200d810} /* (25, 8, 22) {real, imag} */,
  {32'hc1650520, 32'hc0a6bff0} /* (25, 8, 21) {real, imag} */,
  {32'hc1514f4a, 32'h4122fdf0} /* (25, 8, 20) {real, imag} */,
  {32'hc1f60ce2, 32'h4200f814} /* (25, 8, 19) {real, imag} */,
  {32'h41214670, 32'hc20faa91} /* (25, 8, 18) {real, imag} */,
  {32'h41877030, 32'h411cb686} /* (25, 8, 17) {real, imag} */,
  {32'h4103526c, 32'h00000000} /* (25, 8, 16) {real, imag} */,
  {32'h41877030, 32'hc11cb686} /* (25, 8, 15) {real, imag} */,
  {32'h41214670, 32'h420faa91} /* (25, 8, 14) {real, imag} */,
  {32'hc1f60ce2, 32'hc200f814} /* (25, 8, 13) {real, imag} */,
  {32'hc1514f4a, 32'hc122fdf0} /* (25, 8, 12) {real, imag} */,
  {32'hc1650520, 32'h40a6bff0} /* (25, 8, 11) {real, imag} */,
  {32'hc2744fcf, 32'hc200d810} /* (25, 8, 10) {real, imag} */,
  {32'hc2800664, 32'h41bb48fb} /* (25, 8, 9) {real, imag} */,
  {32'hc02618e8, 32'h431cdbf0} /* (25, 8, 8) {real, imag} */,
  {32'hc15ee60e, 32'h429d5b88} /* (25, 8, 7) {real, imag} */,
  {32'hc265d837, 32'h42d7a465} /* (25, 8, 6) {real, imag} */,
  {32'h4201ab4c, 32'h425e7e7e} /* (25, 8, 5) {real, imag} */,
  {32'hc2a8870e, 32'hc194deac} /* (25, 8, 4) {real, imag} */,
  {32'h420200f7, 32'h41abc3e6} /* (25, 8, 3) {real, imag} */,
  {32'h43cbae23, 32'h430589df} /* (25, 8, 2) {real, imag} */,
  {32'hc4c5deb3, 32'hc4569bae} /* (25, 8, 1) {real, imag} */,
  {32'hc4e9802d, 32'h00000000} /* (25, 8, 0) {real, imag} */,
  {32'hc4e3784e, 32'h447daebc} /* (25, 7, 31) {real, imag} */,
  {32'h43c5b2f8, 32'hc2c26112} /* (25, 7, 30) {real, imag} */,
  {32'h42973084, 32'hc192a1dc} /* (25, 7, 29) {real, imag} */,
  {32'hc24e8af0, 32'h4211a301} /* (25, 7, 28) {real, imag} */,
  {32'h435fc39c, 32'hc2cb5593} /* (25, 7, 27) {real, imag} */,
  {32'h421c087c, 32'hc3451a51} /* (25, 7, 26) {real, imag} */,
  {32'hc26635aa, 32'hc2b036bb} /* (25, 7, 25) {real, imag} */,
  {32'hc216d29d, 32'hc32330e9} /* (25, 7, 24) {real, imag} */,
  {32'hc1ed63e7, 32'hc31bbf9c} /* (25, 7, 23) {real, imag} */,
  {32'h4250e09c, 32'h403b18e4} /* (25, 7, 22) {real, imag} */,
  {32'h42e43303, 32'h400d6e60} /* (25, 7, 21) {real, imag} */,
  {32'h4233448f, 32'h420b72fe} /* (25, 7, 20) {real, imag} */,
  {32'h412acb8a, 32'h41bc40a2} /* (25, 7, 19) {real, imag} */,
  {32'hc249bf32, 32'hc1816d5d} /* (25, 7, 18) {real, imag} */,
  {32'h410b87fc, 32'h42498bc4} /* (25, 7, 17) {real, imag} */,
  {32'h407219b0, 32'h00000000} /* (25, 7, 16) {real, imag} */,
  {32'h410b87fc, 32'hc2498bc4} /* (25, 7, 15) {real, imag} */,
  {32'hc249bf32, 32'h41816d5d} /* (25, 7, 14) {real, imag} */,
  {32'h412acb8a, 32'hc1bc40a2} /* (25, 7, 13) {real, imag} */,
  {32'h4233448f, 32'hc20b72fe} /* (25, 7, 12) {real, imag} */,
  {32'h42e43303, 32'hc00d6e60} /* (25, 7, 11) {real, imag} */,
  {32'h4250e09c, 32'hc03b18e4} /* (25, 7, 10) {real, imag} */,
  {32'hc1ed63e7, 32'h431bbf9c} /* (25, 7, 9) {real, imag} */,
  {32'hc216d29d, 32'h432330e9} /* (25, 7, 8) {real, imag} */,
  {32'hc26635aa, 32'h42b036bb} /* (25, 7, 7) {real, imag} */,
  {32'h421c087c, 32'h43451a51} /* (25, 7, 6) {real, imag} */,
  {32'h435fc39c, 32'h42cb5593} /* (25, 7, 5) {real, imag} */,
  {32'hc24e8af0, 32'hc211a301} /* (25, 7, 4) {real, imag} */,
  {32'h42973084, 32'h4192a1dc} /* (25, 7, 3) {real, imag} */,
  {32'h43c5b2f8, 32'h42c26112} /* (25, 7, 2) {real, imag} */,
  {32'hc4e3784e, 32'hc47daebc} /* (25, 7, 1) {real, imag} */,
  {32'hc51c7402, 32'h00000000} /* (25, 7, 0) {real, imag} */,
  {32'hc4eeb672, 32'h449f19ac} /* (25, 6, 31) {real, imag} */,
  {32'h438eabb2, 32'hc361fde2} /* (25, 6, 30) {real, imag} */,
  {32'h42a760df, 32'h401a1018} /* (25, 6, 29) {real, imag} */,
  {32'h4069d918, 32'hc046eb78} /* (25, 6, 28) {real, imag} */,
  {32'h43283f92, 32'h4236c635} /* (25, 6, 27) {real, imag} */,
  {32'h409b52ec, 32'h4249d98e} /* (25, 6, 26) {real, imag} */,
  {32'hc226ce22, 32'hc29a86c2} /* (25, 6, 25) {real, imag} */,
  {32'h405c539c, 32'hc2467c5e} /* (25, 6, 24) {real, imag} */,
  {32'hc1ad2a3f, 32'h4244b5dc} /* (25, 6, 23) {real, imag} */,
  {32'hc1921a72, 32'h423d6f8a} /* (25, 6, 22) {real, imag} */,
  {32'h42cd441a, 32'hc28bdec0} /* (25, 6, 21) {real, imag} */,
  {32'h41c76219, 32'hc1aba3ac} /* (25, 6, 20) {real, imag} */,
  {32'h42909947, 32'hc1c8f45d} /* (25, 6, 19) {real, imag} */,
  {32'h404d09c8, 32'hc1ad2f29} /* (25, 6, 18) {real, imag} */,
  {32'hc23ed11c, 32'h423721cc} /* (25, 6, 17) {real, imag} */,
  {32'h4235dc02, 32'h00000000} /* (25, 6, 16) {real, imag} */,
  {32'hc23ed11c, 32'hc23721cc} /* (25, 6, 15) {real, imag} */,
  {32'h404d09c8, 32'h41ad2f29} /* (25, 6, 14) {real, imag} */,
  {32'h42909947, 32'h41c8f45d} /* (25, 6, 13) {real, imag} */,
  {32'h41c76219, 32'h41aba3ac} /* (25, 6, 12) {real, imag} */,
  {32'h42cd441a, 32'h428bdec0} /* (25, 6, 11) {real, imag} */,
  {32'hc1921a72, 32'hc23d6f8a} /* (25, 6, 10) {real, imag} */,
  {32'hc1ad2a3f, 32'hc244b5dc} /* (25, 6, 9) {real, imag} */,
  {32'h405c539c, 32'h42467c5e} /* (25, 6, 8) {real, imag} */,
  {32'hc226ce22, 32'h429a86c2} /* (25, 6, 7) {real, imag} */,
  {32'h409b52ec, 32'hc249d98e} /* (25, 6, 6) {real, imag} */,
  {32'h43283f92, 32'hc236c635} /* (25, 6, 5) {real, imag} */,
  {32'h4069d918, 32'h4046eb78} /* (25, 6, 4) {real, imag} */,
  {32'h42a760df, 32'hc01a1018} /* (25, 6, 3) {real, imag} */,
  {32'h438eabb2, 32'h4361fde2} /* (25, 6, 2) {real, imag} */,
  {32'hc4eeb672, 32'hc49f19ac} /* (25, 6, 1) {real, imag} */,
  {32'hc521ac05, 32'h00000000} /* (25, 6, 0) {real, imag} */,
  {32'hc4f131eb, 32'h44d0a541} /* (25, 5, 31) {real, imag} */,
  {32'hc1e27130, 32'hc3976bb2} /* (25, 5, 30) {real, imag} */,
  {32'h4077d800, 32'hc1f33cc0} /* (25, 5, 29) {real, imag} */,
  {32'h42aa963d, 32'hc2bdf506} /* (25, 5, 28) {real, imag} */,
  {32'h42ebc65c, 32'h429bde87} /* (25, 5, 27) {real, imag} */,
  {32'h4187a070, 32'h417f1cc0} /* (25, 5, 26) {real, imag} */,
  {32'hc216a22c, 32'hc2b7a825} /* (25, 5, 25) {real, imag} */,
  {32'h420b701d, 32'hc336188a} /* (25, 5, 24) {real, imag} */,
  {32'h41000b34, 32'h413bac4c} /* (25, 5, 23) {real, imag} */,
  {32'h42ac66d9, 32'h41e9f4c2} /* (25, 5, 22) {real, imag} */,
  {32'h427b0e97, 32'h421dd6fe} /* (25, 5, 21) {real, imag} */,
  {32'hc0acfa2c, 32'hc2a78f2d} /* (25, 5, 20) {real, imag} */,
  {32'h410963d7, 32'hc2993b99} /* (25, 5, 19) {real, imag} */,
  {32'h4216fce8, 32'hc2e8b816} /* (25, 5, 18) {real, imag} */,
  {32'h42672e2d, 32'hc277b9da} /* (25, 5, 17) {real, imag} */,
  {32'h42575d11, 32'h00000000} /* (25, 5, 16) {real, imag} */,
  {32'h42672e2d, 32'h4277b9da} /* (25, 5, 15) {real, imag} */,
  {32'h4216fce8, 32'h42e8b816} /* (25, 5, 14) {real, imag} */,
  {32'h410963d7, 32'h42993b99} /* (25, 5, 13) {real, imag} */,
  {32'hc0acfa2c, 32'h42a78f2d} /* (25, 5, 12) {real, imag} */,
  {32'h427b0e97, 32'hc21dd6fe} /* (25, 5, 11) {real, imag} */,
  {32'h42ac66d9, 32'hc1e9f4c2} /* (25, 5, 10) {real, imag} */,
  {32'h41000b34, 32'hc13bac4c} /* (25, 5, 9) {real, imag} */,
  {32'h420b701d, 32'h4336188a} /* (25, 5, 8) {real, imag} */,
  {32'hc216a22c, 32'h42b7a825} /* (25, 5, 7) {real, imag} */,
  {32'h4187a070, 32'hc17f1cc0} /* (25, 5, 6) {real, imag} */,
  {32'h42ebc65c, 32'hc29bde87} /* (25, 5, 5) {real, imag} */,
  {32'h42aa963d, 32'h42bdf506} /* (25, 5, 4) {real, imag} */,
  {32'h4077d800, 32'h41f33cc0} /* (25, 5, 3) {real, imag} */,
  {32'hc1e27130, 32'h43976bb2} /* (25, 5, 2) {real, imag} */,
  {32'hc4f131eb, 32'hc4d0a541} /* (25, 5, 1) {real, imag} */,
  {32'hc5367f94, 32'h00000000} /* (25, 5, 0) {real, imag} */,
  {32'hc4d67225, 32'h450015eb} /* (25, 4, 31) {real, imag} */,
  {32'hc333cd4a, 32'hc386a0c4} /* (25, 4, 30) {real, imag} */,
  {32'h43033608, 32'hc0cf0a50} /* (25, 4, 29) {real, imag} */,
  {32'h42fc3fbc, 32'hc3144d43} /* (25, 4, 28) {real, imag} */,
  {32'h431a9f0f, 32'h4309386d} /* (25, 4, 27) {real, imag} */,
  {32'h41a0118a, 32'hc14871ec} /* (25, 4, 26) {real, imag} */,
  {32'hc2a9a06e, 32'h41bb1912} /* (25, 4, 25) {real, imag} */,
  {32'hc2947c3f, 32'hc238f019} /* (25, 4, 24) {real, imag} */,
  {32'h42be22d4, 32'h423f2f7e} /* (25, 4, 23) {real, imag} */,
  {32'h3f5bc280, 32'hc29b7cf2} /* (25, 4, 22) {real, imag} */,
  {32'h42b36841, 32'hc25f618f} /* (25, 4, 21) {real, imag} */,
  {32'hc0e140b8, 32'h4206e078} /* (25, 4, 20) {real, imag} */,
  {32'hc1ff360c, 32'h429b41be} /* (25, 4, 19) {real, imag} */,
  {32'hc2eb0c5a, 32'h422d0a7c} /* (25, 4, 18) {real, imag} */,
  {32'h416866e8, 32'h41efe3db} /* (25, 4, 17) {real, imag} */,
  {32'h41ade03e, 32'h00000000} /* (25, 4, 16) {real, imag} */,
  {32'h416866e8, 32'hc1efe3db} /* (25, 4, 15) {real, imag} */,
  {32'hc2eb0c5a, 32'hc22d0a7c} /* (25, 4, 14) {real, imag} */,
  {32'hc1ff360c, 32'hc29b41be} /* (25, 4, 13) {real, imag} */,
  {32'hc0e140b8, 32'hc206e078} /* (25, 4, 12) {real, imag} */,
  {32'h42b36841, 32'h425f618f} /* (25, 4, 11) {real, imag} */,
  {32'h3f5bc280, 32'h429b7cf2} /* (25, 4, 10) {real, imag} */,
  {32'h42be22d4, 32'hc23f2f7e} /* (25, 4, 9) {real, imag} */,
  {32'hc2947c3f, 32'h4238f019} /* (25, 4, 8) {real, imag} */,
  {32'hc2a9a06e, 32'hc1bb1912} /* (25, 4, 7) {real, imag} */,
  {32'h41a0118a, 32'h414871ec} /* (25, 4, 6) {real, imag} */,
  {32'h431a9f0f, 32'hc309386d} /* (25, 4, 5) {real, imag} */,
  {32'h42fc3fbc, 32'h43144d43} /* (25, 4, 4) {real, imag} */,
  {32'h43033608, 32'h40cf0a50} /* (25, 4, 3) {real, imag} */,
  {32'hc333cd4a, 32'h4386a0c4} /* (25, 4, 2) {real, imag} */,
  {32'hc4d67225, 32'hc50015eb} /* (25, 4, 1) {real, imag} */,
  {32'hc538b4a2, 32'h00000000} /* (25, 4, 0) {real, imag} */,
  {32'hc4e5f6e4, 32'h450a7f74} /* (25, 3, 31) {real, imag} */,
  {32'hc382f857, 32'hc3b25250} /* (25, 3, 30) {real, imag} */,
  {32'h433f5137, 32'hc296e75c} /* (25, 3, 29) {real, imag} */,
  {32'h4307d455, 32'hc3343270} /* (25, 3, 28) {real, imag} */,
  {32'h43653f7f, 32'hc1ae7124} /* (25, 3, 27) {real, imag} */,
  {32'hc2c376df, 32'h42ab3066} /* (25, 3, 26) {real, imag} */,
  {32'hc2a8a110, 32'hc1fb6c40} /* (25, 3, 25) {real, imag} */,
  {32'hc3437486, 32'hc19d43b8} /* (25, 3, 24) {real, imag} */,
  {32'h42f60d9a, 32'hc1d2a4d4} /* (25, 3, 23) {real, imag} */,
  {32'hc10a3668, 32'hc13e552e} /* (25, 3, 22) {real, imag} */,
  {32'hc18f1cce, 32'hc23a3daf} /* (25, 3, 21) {real, imag} */,
  {32'h4221dcaa, 32'hc2dd5fe5} /* (25, 3, 20) {real, imag} */,
  {32'hbfe2736c, 32'h42a58d88} /* (25, 3, 19) {real, imag} */,
  {32'hc0c932fc, 32'hc1db000c} /* (25, 3, 18) {real, imag} */,
  {32'h42497c6c, 32'h4235188e} /* (25, 3, 17) {real, imag} */,
  {32'hc2a0c2dc, 32'h00000000} /* (25, 3, 16) {real, imag} */,
  {32'h42497c6c, 32'hc235188e} /* (25, 3, 15) {real, imag} */,
  {32'hc0c932fc, 32'h41db000c} /* (25, 3, 14) {real, imag} */,
  {32'hbfe2736c, 32'hc2a58d88} /* (25, 3, 13) {real, imag} */,
  {32'h4221dcaa, 32'h42dd5fe5} /* (25, 3, 12) {real, imag} */,
  {32'hc18f1cce, 32'h423a3daf} /* (25, 3, 11) {real, imag} */,
  {32'hc10a3668, 32'h413e552e} /* (25, 3, 10) {real, imag} */,
  {32'h42f60d9a, 32'h41d2a4d4} /* (25, 3, 9) {real, imag} */,
  {32'hc3437486, 32'h419d43b8} /* (25, 3, 8) {real, imag} */,
  {32'hc2a8a110, 32'h41fb6c40} /* (25, 3, 7) {real, imag} */,
  {32'hc2c376df, 32'hc2ab3066} /* (25, 3, 6) {real, imag} */,
  {32'h43653f7f, 32'h41ae7124} /* (25, 3, 5) {real, imag} */,
  {32'h4307d455, 32'h43343270} /* (25, 3, 4) {real, imag} */,
  {32'h433f5137, 32'h4296e75c} /* (25, 3, 3) {real, imag} */,
  {32'hc382f857, 32'h43b25250} /* (25, 3, 2) {real, imag} */,
  {32'hc4e5f6e4, 32'hc50a7f74} /* (25, 3, 1) {real, imag} */,
  {32'hc5410144, 32'h00000000} /* (25, 3, 0) {real, imag} */,
  {32'hc4ef53e8, 32'h45055565} /* (25, 2, 31) {real, imag} */,
  {32'hc3462532, 32'hc3c65ede} /* (25, 2, 30) {real, imag} */,
  {32'h42ed09d0, 32'h41b81324} /* (25, 2, 29) {real, imag} */,
  {32'h4379712a, 32'hc3437902} /* (25, 2, 28) {real, imag} */,
  {32'h4358bf9c, 32'hc0d9e1b4} /* (25, 2, 27) {real, imag} */,
  {32'h42196829, 32'h421bbbcc} /* (25, 2, 26) {real, imag} */,
  {32'hc2fa8466, 32'h42109b08} /* (25, 2, 25) {real, imag} */,
  {32'hc2e3c692, 32'hc15f2380} /* (25, 2, 24) {real, imag} */,
  {32'hc21e6b4b, 32'hc15967a4} /* (25, 2, 23) {real, imag} */,
  {32'h42f9a972, 32'hc31e97ae} /* (25, 2, 22) {real, imag} */,
  {32'h4287fb57, 32'h4240e662} /* (25, 2, 21) {real, imag} */,
  {32'hc182c281, 32'h427c336c} /* (25, 2, 20) {real, imag} */,
  {32'hc24e7b53, 32'hc2b067c7} /* (25, 2, 19) {real, imag} */,
  {32'hc188f25e, 32'hc101bfd0} /* (25, 2, 18) {real, imag} */,
  {32'h41c70b97, 32'hc1832c2f} /* (25, 2, 17) {real, imag} */,
  {32'hc2743cd0, 32'h00000000} /* (25, 2, 16) {real, imag} */,
  {32'h41c70b97, 32'h41832c2f} /* (25, 2, 15) {real, imag} */,
  {32'hc188f25e, 32'h4101bfd0} /* (25, 2, 14) {real, imag} */,
  {32'hc24e7b53, 32'h42b067c7} /* (25, 2, 13) {real, imag} */,
  {32'hc182c281, 32'hc27c336c} /* (25, 2, 12) {real, imag} */,
  {32'h4287fb57, 32'hc240e662} /* (25, 2, 11) {real, imag} */,
  {32'h42f9a972, 32'h431e97ae} /* (25, 2, 10) {real, imag} */,
  {32'hc21e6b4b, 32'h415967a4} /* (25, 2, 9) {real, imag} */,
  {32'hc2e3c692, 32'h415f2380} /* (25, 2, 8) {real, imag} */,
  {32'hc2fa8466, 32'hc2109b08} /* (25, 2, 7) {real, imag} */,
  {32'h42196829, 32'hc21bbbcc} /* (25, 2, 6) {real, imag} */,
  {32'h4358bf9c, 32'h40d9e1b4} /* (25, 2, 5) {real, imag} */,
  {32'h4379712a, 32'h43437902} /* (25, 2, 4) {real, imag} */,
  {32'h42ed09d0, 32'hc1b81324} /* (25, 2, 3) {real, imag} */,
  {32'hc3462532, 32'h43c65ede} /* (25, 2, 2) {real, imag} */,
  {32'hc4ef53e8, 32'hc5055565} /* (25, 2, 1) {real, imag} */,
  {32'hc53aac66, 32'h00000000} /* (25, 2, 0) {real, imag} */,
  {32'hc4e4754a, 32'h44eb03be} /* (25, 1, 31) {real, imag} */,
  {32'hc2ec5592, 32'hc38d8dc2} /* (25, 1, 30) {real, imag} */,
  {32'h433f3ac8, 32'h418cc148} /* (25, 1, 29) {real, imag} */,
  {32'h433c6478, 32'hc2af5062} /* (25, 1, 28) {real, imag} */,
  {32'h42981e3e, 32'h419d3295} /* (25, 1, 27) {real, imag} */,
  {32'hc264dff7, 32'hc27d0008} /* (25, 1, 26) {real, imag} */,
  {32'h425bf5d2, 32'h42d18242} /* (25, 1, 25) {real, imag} */,
  {32'hc2a9907f, 32'hc2966ddc} /* (25, 1, 24) {real, imag} */,
  {32'h4293138e, 32'h42c3de0b} /* (25, 1, 23) {real, imag} */,
  {32'hc23da8d5, 32'hc14fd245} /* (25, 1, 22) {real, imag} */,
  {32'h429f2295, 32'hc2a34f16} /* (25, 1, 21) {real, imag} */,
  {32'hc1873248, 32'h418c8ea0} /* (25, 1, 20) {real, imag} */,
  {32'h42aad471, 32'hc213b165} /* (25, 1, 19) {real, imag} */,
  {32'hc29606cd, 32'hc2a3de5d} /* (25, 1, 18) {real, imag} */,
  {32'hc2d61a1e, 32'hc09c69fd} /* (25, 1, 17) {real, imag} */,
  {32'h40ab7418, 32'h00000000} /* (25, 1, 16) {real, imag} */,
  {32'hc2d61a1e, 32'h409c69fd} /* (25, 1, 15) {real, imag} */,
  {32'hc29606cd, 32'h42a3de5d} /* (25, 1, 14) {real, imag} */,
  {32'h42aad471, 32'h4213b165} /* (25, 1, 13) {real, imag} */,
  {32'hc1873248, 32'hc18c8ea0} /* (25, 1, 12) {real, imag} */,
  {32'h429f2295, 32'h42a34f16} /* (25, 1, 11) {real, imag} */,
  {32'hc23da8d5, 32'h414fd245} /* (25, 1, 10) {real, imag} */,
  {32'h4293138e, 32'hc2c3de0b} /* (25, 1, 9) {real, imag} */,
  {32'hc2a9907f, 32'h42966ddc} /* (25, 1, 8) {real, imag} */,
  {32'h425bf5d2, 32'hc2d18242} /* (25, 1, 7) {real, imag} */,
  {32'hc264dff7, 32'h427d0008} /* (25, 1, 6) {real, imag} */,
  {32'h42981e3e, 32'hc19d3295} /* (25, 1, 5) {real, imag} */,
  {32'h433c6478, 32'h42af5062} /* (25, 1, 4) {real, imag} */,
  {32'h433f3ac8, 32'hc18cc148} /* (25, 1, 3) {real, imag} */,
  {32'hc2ec5592, 32'h438d8dc2} /* (25, 1, 2) {real, imag} */,
  {32'hc4e4754a, 32'hc4eb03be} /* (25, 1, 1) {real, imag} */,
  {32'hc543edb7, 32'h00000000} /* (25, 1, 0) {real, imag} */,
  {32'hc4ee5faf, 32'h44b34140} /* (25, 0, 31) {real, imag} */,
  {32'h42849714, 32'hc32c8d2d} /* (25, 0, 30) {real, imag} */,
  {32'h42d944ce, 32'hc28f699c} /* (25, 0, 29) {real, imag} */,
  {32'h424c616f, 32'hc2cbb264} /* (25, 0, 28) {real, imag} */,
  {32'h42c7db05, 32'hc2ae9e5c} /* (25, 0, 27) {real, imag} */,
  {32'hc1de39ce, 32'hc1f9812c} /* (25, 0, 26) {real, imag} */,
  {32'h40a3b3a2, 32'h41e20e5e} /* (25, 0, 25) {real, imag} */,
  {32'h426c90ec, 32'hc232bdd1} /* (25, 0, 24) {real, imag} */,
  {32'h4225d5dc, 32'h40934a68} /* (25, 0, 23) {real, imag} */,
  {32'h42430a5e, 32'h3fe9b800} /* (25, 0, 22) {real, imag} */,
  {32'h40f91300, 32'h41ed8f0e} /* (25, 0, 21) {real, imag} */,
  {32'h41fe72a5, 32'h4150f398} /* (25, 0, 20) {real, imag} */,
  {32'h4216a5e4, 32'h4229477a} /* (25, 0, 19) {real, imag} */,
  {32'h42373990, 32'h41286952} /* (25, 0, 18) {real, imag} */,
  {32'hc11fe97c, 32'hc1b564d8} /* (25, 0, 17) {real, imag} */,
  {32'h410a4638, 32'h00000000} /* (25, 0, 16) {real, imag} */,
  {32'hc11fe97c, 32'h41b564d8} /* (25, 0, 15) {real, imag} */,
  {32'h42373990, 32'hc1286952} /* (25, 0, 14) {real, imag} */,
  {32'h4216a5e4, 32'hc229477a} /* (25, 0, 13) {real, imag} */,
  {32'h41fe72a5, 32'hc150f398} /* (25, 0, 12) {real, imag} */,
  {32'h40f91300, 32'hc1ed8f0e} /* (25, 0, 11) {real, imag} */,
  {32'h42430a5e, 32'hbfe9b800} /* (25, 0, 10) {real, imag} */,
  {32'h4225d5dc, 32'hc0934a68} /* (25, 0, 9) {real, imag} */,
  {32'h426c90ec, 32'h4232bdd1} /* (25, 0, 8) {real, imag} */,
  {32'h40a3b3a2, 32'hc1e20e5e} /* (25, 0, 7) {real, imag} */,
  {32'hc1de39ce, 32'h41f9812c} /* (25, 0, 6) {real, imag} */,
  {32'h42c7db05, 32'h42ae9e5c} /* (25, 0, 5) {real, imag} */,
  {32'h424c616f, 32'h42cbb264} /* (25, 0, 4) {real, imag} */,
  {32'h42d944ce, 32'h428f699c} /* (25, 0, 3) {real, imag} */,
  {32'h42849714, 32'h432c8d2d} /* (25, 0, 2) {real, imag} */,
  {32'hc4ee5faf, 32'hc4b34140} /* (25, 0, 1) {real, imag} */,
  {32'hc53f26a0, 32'h00000000} /* (25, 0, 0) {real, imag} */,
  {32'hc53fc377, 32'h44d32d0c} /* (24, 31, 31) {real, imag} */,
  {32'h4414a04e, 32'hc31e99e5} /* (24, 31, 30) {real, imag} */,
  {32'h429f7337, 32'hbe982ea0} /* (24, 31, 29) {real, imag} */,
  {32'hc214feee, 32'h40aa92a0} /* (24, 31, 28) {real, imag} */,
  {32'h43306db6, 32'hc21f25e4} /* (24, 31, 27) {real, imag} */,
  {32'hc285f85e, 32'hc1925e98} /* (24, 31, 26) {real, imag} */,
  {32'hc2442882, 32'h410d6210} /* (24, 31, 25) {real, imag} */,
  {32'h427eb2e6, 32'hc2994b8e} /* (24, 31, 24) {real, imag} */,
  {32'h41c1bb11, 32'h41c563f5} /* (24, 31, 23) {real, imag} */,
  {32'h42b8033a, 32'hc1c8be61} /* (24, 31, 22) {real, imag} */,
  {32'h416771cb, 32'hc254c01e} /* (24, 31, 21) {real, imag} */,
  {32'hc222fa68, 32'h3fd6c000} /* (24, 31, 20) {real, imag} */,
  {32'hc2b51c7a, 32'hc212b79f} /* (24, 31, 19) {real, imag} */,
  {32'h4281f771, 32'h41ceadaa} /* (24, 31, 18) {real, imag} */,
  {32'h41f35b58, 32'h42307912} /* (24, 31, 17) {real, imag} */,
  {32'hc271e948, 32'h00000000} /* (24, 31, 16) {real, imag} */,
  {32'h41f35b58, 32'hc2307912} /* (24, 31, 15) {real, imag} */,
  {32'h4281f771, 32'hc1ceadaa} /* (24, 31, 14) {real, imag} */,
  {32'hc2b51c7a, 32'h4212b79f} /* (24, 31, 13) {real, imag} */,
  {32'hc222fa68, 32'hbfd6c000} /* (24, 31, 12) {real, imag} */,
  {32'h416771cb, 32'h4254c01e} /* (24, 31, 11) {real, imag} */,
  {32'h42b8033a, 32'h41c8be61} /* (24, 31, 10) {real, imag} */,
  {32'h41c1bb11, 32'hc1c563f5} /* (24, 31, 9) {real, imag} */,
  {32'h427eb2e6, 32'h42994b8e} /* (24, 31, 8) {real, imag} */,
  {32'hc2442882, 32'hc10d6210} /* (24, 31, 7) {real, imag} */,
  {32'hc285f85e, 32'h41925e98} /* (24, 31, 6) {real, imag} */,
  {32'h43306db6, 32'h421f25e4} /* (24, 31, 5) {real, imag} */,
  {32'hc214feee, 32'hc0aa92a0} /* (24, 31, 4) {real, imag} */,
  {32'h429f7337, 32'h3e982ea0} /* (24, 31, 3) {real, imag} */,
  {32'h4414a04e, 32'h431e99e5} /* (24, 31, 2) {real, imag} */,
  {32'hc53fc377, 32'hc4d32d0c} /* (24, 31, 1) {real, imag} */,
  {32'hc58502ae, 32'h00000000} /* (24, 31, 0) {real, imag} */,
  {32'hc55bd0bd, 32'h44ae15cc} /* (24, 30, 31) {real, imag} */,
  {32'h4470354b, 32'hc354e104} /* (24, 30, 30) {real, imag} */,
  {32'h42c57a62, 32'hc1de4250} /* (24, 30, 29) {real, imag} */,
  {32'hc2c3dd1c, 32'h42ec1666} /* (24, 30, 28) {real, imag} */,
  {32'h43255736, 32'hc2fe7f18} /* (24, 30, 27) {real, imag} */,
  {32'h41468c2c, 32'h406a0898} /* (24, 30, 26) {real, imag} */,
  {32'hc216560d, 32'h4289df1b} /* (24, 30, 25) {real, imag} */,
  {32'h42db5479, 32'hc2601416} /* (24, 30, 24) {real, imag} */,
  {32'h41a2099d, 32'hc18a4342} /* (24, 30, 23) {real, imag} */,
  {32'hc22e486c, 32'h42ebd3e8} /* (24, 30, 22) {real, imag} */,
  {32'h42cc9068, 32'hc2858edc} /* (24, 30, 21) {real, imag} */,
  {32'hc2774e6c, 32'hc21a9b30} /* (24, 30, 20) {real, imag} */,
  {32'hc2d578e5, 32'hc2068806} /* (24, 30, 19) {real, imag} */,
  {32'h4263c3c7, 32'hc1eadc94} /* (24, 30, 18) {real, imag} */,
  {32'hc0cb6ba8, 32'h4268b330} /* (24, 30, 17) {real, imag} */,
  {32'h41460f00, 32'h00000000} /* (24, 30, 16) {real, imag} */,
  {32'hc0cb6ba8, 32'hc268b330} /* (24, 30, 15) {real, imag} */,
  {32'h4263c3c7, 32'h41eadc94} /* (24, 30, 14) {real, imag} */,
  {32'hc2d578e5, 32'h42068806} /* (24, 30, 13) {real, imag} */,
  {32'hc2774e6c, 32'h421a9b30} /* (24, 30, 12) {real, imag} */,
  {32'h42cc9068, 32'h42858edc} /* (24, 30, 11) {real, imag} */,
  {32'hc22e486c, 32'hc2ebd3e8} /* (24, 30, 10) {real, imag} */,
  {32'h41a2099d, 32'h418a4342} /* (24, 30, 9) {real, imag} */,
  {32'h42db5479, 32'h42601416} /* (24, 30, 8) {real, imag} */,
  {32'hc216560d, 32'hc289df1b} /* (24, 30, 7) {real, imag} */,
  {32'h41468c2c, 32'hc06a0898} /* (24, 30, 6) {real, imag} */,
  {32'h43255736, 32'h42fe7f18} /* (24, 30, 5) {real, imag} */,
  {32'hc2c3dd1c, 32'hc2ec1666} /* (24, 30, 4) {real, imag} */,
  {32'h42c57a62, 32'h41de4250} /* (24, 30, 3) {real, imag} */,
  {32'h4470354b, 32'h4354e104} /* (24, 30, 2) {real, imag} */,
  {32'hc55bd0bd, 32'hc4ae15cc} /* (24, 30, 1) {real, imag} */,
  {32'hc585ed5b, 32'h00000000} /* (24, 30, 0) {real, imag} */,
  {32'hc56818bc, 32'h449ceaea} /* (24, 29, 31) {real, imag} */,
  {32'h4480848d, 32'hc2fa18dc} /* (24, 29, 30) {real, imag} */,
  {32'h42384fc8, 32'h412a08f8} /* (24, 29, 29) {real, imag} */,
  {32'hc366caf7, 32'h4286c01e} /* (24, 29, 28) {real, imag} */,
  {32'h42b88df0, 32'hc3107f8a} /* (24, 29, 27) {real, imag} */,
  {32'h43103b84, 32'hc1af3726} /* (24, 29, 26) {real, imag} */,
  {32'h430e0da0, 32'h41d7b064} /* (24, 29, 25) {real, imag} */,
  {32'h42d0c745, 32'h40b220b8} /* (24, 29, 24) {real, imag} */,
  {32'hc25e33f3, 32'hc19917b5} /* (24, 29, 23) {real, imag} */,
  {32'hc22b9519, 32'h413e5978} /* (24, 29, 22) {real, imag} */,
  {32'h42543325, 32'h41531621} /* (24, 29, 21) {real, imag} */,
  {32'hc2b71993, 32'hc1b577e5} /* (24, 29, 20) {real, imag} */,
  {32'hc2984f11, 32'hc22ed8b4} /* (24, 29, 19) {real, imag} */,
  {32'hc1fd19d8, 32'hc21bc49d} /* (24, 29, 18) {real, imag} */,
  {32'hc15335f2, 32'hc245adba} /* (24, 29, 17) {real, imag} */,
  {32'h42e0d8df, 32'h00000000} /* (24, 29, 16) {real, imag} */,
  {32'hc15335f2, 32'h4245adba} /* (24, 29, 15) {real, imag} */,
  {32'hc1fd19d8, 32'h421bc49d} /* (24, 29, 14) {real, imag} */,
  {32'hc2984f11, 32'h422ed8b4} /* (24, 29, 13) {real, imag} */,
  {32'hc2b71993, 32'h41b577e5} /* (24, 29, 12) {real, imag} */,
  {32'h42543325, 32'hc1531621} /* (24, 29, 11) {real, imag} */,
  {32'hc22b9519, 32'hc13e5978} /* (24, 29, 10) {real, imag} */,
  {32'hc25e33f3, 32'h419917b5} /* (24, 29, 9) {real, imag} */,
  {32'h42d0c745, 32'hc0b220b8} /* (24, 29, 8) {real, imag} */,
  {32'h430e0da0, 32'hc1d7b064} /* (24, 29, 7) {real, imag} */,
  {32'h43103b84, 32'h41af3726} /* (24, 29, 6) {real, imag} */,
  {32'h42b88df0, 32'h43107f8a} /* (24, 29, 5) {real, imag} */,
  {32'hc366caf7, 32'hc286c01e} /* (24, 29, 4) {real, imag} */,
  {32'h42384fc8, 32'hc12a08f8} /* (24, 29, 3) {real, imag} */,
  {32'h4480848d, 32'h42fa18dc} /* (24, 29, 2) {real, imag} */,
  {32'hc56818bc, 32'hc49ceaea} /* (24, 29, 1) {real, imag} */,
  {32'hc5888115, 32'h00000000} /* (24, 29, 0) {real, imag} */,
  {32'hc575f335, 32'h448a97c2} /* (24, 28, 31) {real, imag} */,
  {32'h449414e1, 32'hc32e60a8} /* (24, 28, 30) {real, imag} */,
  {32'hc2e7b16e, 32'hc229454c} /* (24, 28, 29) {real, imag} */,
  {32'hc310fe04, 32'h42c53e8a} /* (24, 28, 28) {real, imag} */,
  {32'h431b55f1, 32'hc35d9435} /* (24, 28, 27) {real, imag} */,
  {32'h42a0f53e, 32'h421aca98} /* (24, 28, 26) {real, imag} */,
  {32'hc1f76e2e, 32'h4304b31c} /* (24, 28, 25) {real, imag} */,
  {32'h42f963b2, 32'hc2e7850e} /* (24, 28, 24) {real, imag} */,
  {32'hc21bd78e, 32'h408a9b64} /* (24, 28, 23) {real, imag} */,
  {32'hc28be113, 32'hc2cc70f8} /* (24, 28, 22) {real, imag} */,
  {32'hc292c13a, 32'hc302b109} /* (24, 28, 21) {real, imag} */,
  {32'h417fc4b2, 32'h420a3f8b} /* (24, 28, 20) {real, imag} */,
  {32'h4159c22c, 32'h4256ab72} /* (24, 28, 19) {real, imag} */,
  {32'h419f5099, 32'hc29ca680} /* (24, 28, 18) {real, imag} */,
  {32'h4100fbe0, 32'hc1578f62} /* (24, 28, 17) {real, imag} */,
  {32'hc237bea6, 32'h00000000} /* (24, 28, 16) {real, imag} */,
  {32'h4100fbe0, 32'h41578f62} /* (24, 28, 15) {real, imag} */,
  {32'h419f5099, 32'h429ca680} /* (24, 28, 14) {real, imag} */,
  {32'h4159c22c, 32'hc256ab72} /* (24, 28, 13) {real, imag} */,
  {32'h417fc4b2, 32'hc20a3f8b} /* (24, 28, 12) {real, imag} */,
  {32'hc292c13a, 32'h4302b109} /* (24, 28, 11) {real, imag} */,
  {32'hc28be113, 32'h42cc70f8} /* (24, 28, 10) {real, imag} */,
  {32'hc21bd78e, 32'hc08a9b64} /* (24, 28, 9) {real, imag} */,
  {32'h42f963b2, 32'h42e7850e} /* (24, 28, 8) {real, imag} */,
  {32'hc1f76e2e, 32'hc304b31c} /* (24, 28, 7) {real, imag} */,
  {32'h42a0f53e, 32'hc21aca98} /* (24, 28, 6) {real, imag} */,
  {32'h431b55f1, 32'h435d9435} /* (24, 28, 5) {real, imag} */,
  {32'hc310fe04, 32'hc2c53e8a} /* (24, 28, 4) {real, imag} */,
  {32'hc2e7b16e, 32'h4229454c} /* (24, 28, 3) {real, imag} */,
  {32'h449414e1, 32'h432e60a8} /* (24, 28, 2) {real, imag} */,
  {32'hc575f335, 32'hc48a97c2} /* (24, 28, 1) {real, imag} */,
  {32'hc58ec3c9, 32'h00000000} /* (24, 28, 0) {real, imag} */,
  {32'hc570f256, 32'h447a9168} /* (24, 27, 31) {real, imag} */,
  {32'h449e3028, 32'hc3494f11} /* (24, 27, 30) {real, imag} */,
  {32'h422c2614, 32'hc3527e47} /* (24, 27, 29) {real, imag} */,
  {32'hc32955a0, 32'hc039b320} /* (24, 27, 28) {real, imag} */,
  {32'h431d3f60, 32'hc33f122e} /* (24, 27, 27) {real, imag} */,
  {32'h4207023b, 32'h438ac11e} /* (24, 27, 26) {real, imag} */,
  {32'h413d6f8e, 32'h42483658} /* (24, 27, 25) {real, imag} */,
  {32'h42a1fa50, 32'hc30040ca} /* (24, 27, 24) {real, imag} */,
  {32'h4283b3c7, 32'hc1af78a2} /* (24, 27, 23) {real, imag} */,
  {32'hc29b919e, 32'hc28337ea} /* (24, 27, 22) {real, imag} */,
  {32'hc29d701d, 32'h41f5c960} /* (24, 27, 21) {real, imag} */,
  {32'h424093be, 32'h424d49ca} /* (24, 27, 20) {real, imag} */,
  {32'h4281bb18, 32'h41dc12de} /* (24, 27, 19) {real, imag} */,
  {32'h42833435, 32'hc290782c} /* (24, 27, 18) {real, imag} */,
  {32'h41619245, 32'h422a39e6} /* (24, 27, 17) {real, imag} */,
  {32'hc2587241, 32'h00000000} /* (24, 27, 16) {real, imag} */,
  {32'h41619245, 32'hc22a39e6} /* (24, 27, 15) {real, imag} */,
  {32'h42833435, 32'h4290782c} /* (24, 27, 14) {real, imag} */,
  {32'h4281bb18, 32'hc1dc12de} /* (24, 27, 13) {real, imag} */,
  {32'h424093be, 32'hc24d49ca} /* (24, 27, 12) {real, imag} */,
  {32'hc29d701d, 32'hc1f5c960} /* (24, 27, 11) {real, imag} */,
  {32'hc29b919e, 32'h428337ea} /* (24, 27, 10) {real, imag} */,
  {32'h4283b3c7, 32'h41af78a2} /* (24, 27, 9) {real, imag} */,
  {32'h42a1fa50, 32'h430040ca} /* (24, 27, 8) {real, imag} */,
  {32'h413d6f8e, 32'hc2483658} /* (24, 27, 7) {real, imag} */,
  {32'h4207023b, 32'hc38ac11e} /* (24, 27, 6) {real, imag} */,
  {32'h431d3f60, 32'h433f122e} /* (24, 27, 5) {real, imag} */,
  {32'hc32955a0, 32'h4039b320} /* (24, 27, 4) {real, imag} */,
  {32'h422c2614, 32'h43527e47} /* (24, 27, 3) {real, imag} */,
  {32'h449e3028, 32'h43494f11} /* (24, 27, 2) {real, imag} */,
  {32'hc570f256, 32'hc47a9168} /* (24, 27, 1) {real, imag} */,
  {32'hc58ad12b, 32'h00000000} /* (24, 27, 0) {real, imag} */,
  {32'hc565d2ab, 32'h444b37fc} /* (24, 26, 31) {real, imag} */,
  {32'h44a78be2, 32'hc20d8770} /* (24, 26, 30) {real, imag} */,
  {32'h41e2609e, 32'hc2e22750} /* (24, 26, 29) {real, imag} */,
  {32'hc28aea6c, 32'hc27fa1a5} /* (24, 26, 28) {real, imag} */,
  {32'h4312ae7c, 32'hc2a70042} /* (24, 26, 27) {real, imag} */,
  {32'hc26f4ca4, 32'h432a4e00} /* (24, 26, 26) {real, imag} */,
  {32'h427560c2, 32'h4223e65f} /* (24, 26, 25) {real, imag} */,
  {32'h42f82334, 32'hc24865fe} /* (24, 26, 24) {real, imag} */,
  {32'hc14ced4a, 32'h42503c18} /* (24, 26, 23) {real, imag} */,
  {32'hc226f18c, 32'hc267ae35} /* (24, 26, 22) {real, imag} */,
  {32'hc214faa2, 32'hc230b932} /* (24, 26, 21) {real, imag} */,
  {32'hc22e0034, 32'h4227fabe} /* (24, 26, 20) {real, imag} */,
  {32'h414ed562, 32'hc1e1103b} /* (24, 26, 19) {real, imag} */,
  {32'hc033fe40, 32'hc1deb6a6} /* (24, 26, 18) {real, imag} */,
  {32'hc2595fb2, 32'hc1cb814c} /* (24, 26, 17) {real, imag} */,
  {32'h42a8c0d6, 32'h00000000} /* (24, 26, 16) {real, imag} */,
  {32'hc2595fb2, 32'h41cb814c} /* (24, 26, 15) {real, imag} */,
  {32'hc033fe40, 32'h41deb6a6} /* (24, 26, 14) {real, imag} */,
  {32'h414ed562, 32'h41e1103b} /* (24, 26, 13) {real, imag} */,
  {32'hc22e0034, 32'hc227fabe} /* (24, 26, 12) {real, imag} */,
  {32'hc214faa2, 32'h4230b932} /* (24, 26, 11) {real, imag} */,
  {32'hc226f18c, 32'h4267ae35} /* (24, 26, 10) {real, imag} */,
  {32'hc14ced4a, 32'hc2503c18} /* (24, 26, 9) {real, imag} */,
  {32'h42f82334, 32'h424865fe} /* (24, 26, 8) {real, imag} */,
  {32'h427560c2, 32'hc223e65f} /* (24, 26, 7) {real, imag} */,
  {32'hc26f4ca4, 32'hc32a4e00} /* (24, 26, 6) {real, imag} */,
  {32'h4312ae7c, 32'h42a70042} /* (24, 26, 5) {real, imag} */,
  {32'hc28aea6c, 32'h427fa1a5} /* (24, 26, 4) {real, imag} */,
  {32'h41e2609e, 32'h42e22750} /* (24, 26, 3) {real, imag} */,
  {32'h44a78be2, 32'h420d8770} /* (24, 26, 2) {real, imag} */,
  {32'hc565d2ab, 32'hc44b37fc} /* (24, 26, 1) {real, imag} */,
  {32'hc5830d28, 32'h00000000} /* (24, 26, 0) {real, imag} */,
  {32'hc5619377, 32'h44014af7} /* (24, 25, 31) {real, imag} */,
  {32'h449cd62f, 32'h42ab27b7} /* (24, 25, 30) {real, imag} */,
  {32'h41ec7d36, 32'h4094e804} /* (24, 25, 29) {real, imag} */,
  {32'hc2ac581b, 32'hc107c196} /* (24, 25, 28) {real, imag} */,
  {32'h43762912, 32'hc13f8434} /* (24, 25, 27) {real, imag} */,
  {32'h418370ae, 32'h42924c66} /* (24, 25, 26) {real, imag} */,
  {32'h422db566, 32'h42022314} /* (24, 25, 25) {real, imag} */,
  {32'hc2b59be1, 32'hc2272bd2} /* (24, 25, 24) {real, imag} */,
  {32'hc299ccbc, 32'hc3310993} /* (24, 25, 23) {real, imag} */,
  {32'hc27e2189, 32'hc0897450} /* (24, 25, 22) {real, imag} */,
  {32'h41bc76bc, 32'hc2bfd223} /* (24, 25, 21) {real, imag} */,
  {32'hc28f6c66, 32'h41bd69c9} /* (24, 25, 20) {real, imag} */,
  {32'hc1dce381, 32'hc1e3bcd6} /* (24, 25, 19) {real, imag} */,
  {32'hc2afbcd8, 32'h42b7c5a2} /* (24, 25, 18) {real, imag} */,
  {32'h41d5f269, 32'h41f203f0} /* (24, 25, 17) {real, imag} */,
  {32'h41a8ac09, 32'h00000000} /* (24, 25, 16) {real, imag} */,
  {32'h41d5f269, 32'hc1f203f0} /* (24, 25, 15) {real, imag} */,
  {32'hc2afbcd8, 32'hc2b7c5a2} /* (24, 25, 14) {real, imag} */,
  {32'hc1dce381, 32'h41e3bcd6} /* (24, 25, 13) {real, imag} */,
  {32'hc28f6c66, 32'hc1bd69c9} /* (24, 25, 12) {real, imag} */,
  {32'h41bc76bc, 32'h42bfd223} /* (24, 25, 11) {real, imag} */,
  {32'hc27e2189, 32'h40897450} /* (24, 25, 10) {real, imag} */,
  {32'hc299ccbc, 32'h43310993} /* (24, 25, 9) {real, imag} */,
  {32'hc2b59be1, 32'h42272bd2} /* (24, 25, 8) {real, imag} */,
  {32'h422db566, 32'hc2022314} /* (24, 25, 7) {real, imag} */,
  {32'h418370ae, 32'hc2924c66} /* (24, 25, 6) {real, imag} */,
  {32'h43762912, 32'h413f8434} /* (24, 25, 5) {real, imag} */,
  {32'hc2ac581b, 32'h4107c196} /* (24, 25, 4) {real, imag} */,
  {32'h41ec7d36, 32'hc094e804} /* (24, 25, 3) {real, imag} */,
  {32'h449cd62f, 32'hc2ab27b7} /* (24, 25, 2) {real, imag} */,
  {32'hc5619377, 32'hc4014af7} /* (24, 25, 1) {real, imag} */,
  {32'hc576c0c2, 32'h00000000} /* (24, 25, 0) {real, imag} */,
  {32'hc544b1d2, 32'h43e29bf4} /* (24, 24, 31) {real, imag} */,
  {32'h44939cad, 32'hc2af7668} /* (24, 24, 30) {real, imag} */,
  {32'hc2f8eaaa, 32'hc19ccfc6} /* (24, 24, 29) {real, imag} */,
  {32'hc2c7cebe, 32'hc2a1da5e} /* (24, 24, 28) {real, imag} */,
  {32'h43318e06, 32'hc232fa8c} /* (24, 24, 27) {real, imag} */,
  {32'h42f1fd46, 32'h4107fb18} /* (24, 24, 26) {real, imag} */,
  {32'h42344734, 32'h423a8796} /* (24, 24, 25) {real, imag} */,
  {32'hc242d02a, 32'hc1eebf8f} /* (24, 24, 24) {real, imag} */,
  {32'hc268a302, 32'h3f9e36e8} /* (24, 24, 23) {real, imag} */,
  {32'hc1c85b3a, 32'h42a856ee} /* (24, 24, 22) {real, imag} */,
  {32'hc2769ddf, 32'hc220c7ea} /* (24, 24, 21) {real, imag} */,
  {32'hc17dbb54, 32'h426022c7} /* (24, 24, 20) {real, imag} */,
  {32'hbe8bd160, 32'hc2826fdd} /* (24, 24, 19) {real, imag} */,
  {32'h3f8a8980, 32'hc308281c} /* (24, 24, 18) {real, imag} */,
  {32'hc16b7b3c, 32'h41a6e456} /* (24, 24, 17) {real, imag} */,
  {32'hc18ad264, 32'h00000000} /* (24, 24, 16) {real, imag} */,
  {32'hc16b7b3c, 32'hc1a6e456} /* (24, 24, 15) {real, imag} */,
  {32'h3f8a8980, 32'h4308281c} /* (24, 24, 14) {real, imag} */,
  {32'hbe8bd160, 32'h42826fdd} /* (24, 24, 13) {real, imag} */,
  {32'hc17dbb54, 32'hc26022c7} /* (24, 24, 12) {real, imag} */,
  {32'hc2769ddf, 32'h4220c7ea} /* (24, 24, 11) {real, imag} */,
  {32'hc1c85b3a, 32'hc2a856ee} /* (24, 24, 10) {real, imag} */,
  {32'hc268a302, 32'hbf9e36e8} /* (24, 24, 9) {real, imag} */,
  {32'hc242d02a, 32'h41eebf8f} /* (24, 24, 8) {real, imag} */,
  {32'h42344734, 32'hc23a8796} /* (24, 24, 7) {real, imag} */,
  {32'h42f1fd46, 32'hc107fb18} /* (24, 24, 6) {real, imag} */,
  {32'h43318e06, 32'h4232fa8c} /* (24, 24, 5) {real, imag} */,
  {32'hc2c7cebe, 32'h42a1da5e} /* (24, 24, 4) {real, imag} */,
  {32'hc2f8eaaa, 32'h419ccfc6} /* (24, 24, 3) {real, imag} */,
  {32'h44939cad, 32'h42af7668} /* (24, 24, 2) {real, imag} */,
  {32'hc544b1d2, 32'hc3e29bf4} /* (24, 24, 1) {real, imag} */,
  {32'hc554edb6, 32'h00000000} /* (24, 24, 0) {real, imag} */,
  {32'hc529e172, 32'h43bbc3f2} /* (24, 23, 31) {real, imag} */,
  {32'h44850fde, 32'hc3418478} /* (24, 23, 30) {real, imag} */,
  {32'hc2bb865c, 32'h419b8ca6} /* (24, 23, 29) {real, imag} */,
  {32'hc326d0c5, 32'h41ce6c5a} /* (24, 23, 28) {real, imag} */,
  {32'h4304d756, 32'hc2c1fc15} /* (24, 23, 27) {real, imag} */,
  {32'hc2d13736, 32'hc304b6c8} /* (24, 23, 26) {real, imag} */,
  {32'hc14afbc0, 32'hc1aac09f} /* (24, 23, 25) {real, imag} */,
  {32'h41ffc040, 32'hc28f4603} /* (24, 23, 24) {real, imag} */,
  {32'h42dcf3c2, 32'hc3063a6d} /* (24, 23, 23) {real, imag} */,
  {32'hc188e122, 32'hc22fee56} /* (24, 23, 22) {real, imag} */,
  {32'h42db27f0, 32'hc1e240f0} /* (24, 23, 21) {real, imag} */,
  {32'hc25445f5, 32'h426ee038} /* (24, 23, 20) {real, imag} */,
  {32'hc25c12f1, 32'h41b8c9f4} /* (24, 23, 19) {real, imag} */,
  {32'h420dfab8, 32'hc1a81064} /* (24, 23, 18) {real, imag} */,
  {32'h4050eeae, 32'hc1b181b3} /* (24, 23, 17) {real, imag} */,
  {32'h4263895d, 32'h00000000} /* (24, 23, 16) {real, imag} */,
  {32'h4050eeae, 32'h41b181b3} /* (24, 23, 15) {real, imag} */,
  {32'h420dfab8, 32'h41a81064} /* (24, 23, 14) {real, imag} */,
  {32'hc25c12f1, 32'hc1b8c9f4} /* (24, 23, 13) {real, imag} */,
  {32'hc25445f5, 32'hc26ee038} /* (24, 23, 12) {real, imag} */,
  {32'h42db27f0, 32'h41e240f0} /* (24, 23, 11) {real, imag} */,
  {32'hc188e122, 32'h422fee56} /* (24, 23, 10) {real, imag} */,
  {32'h42dcf3c2, 32'h43063a6d} /* (24, 23, 9) {real, imag} */,
  {32'h41ffc040, 32'h428f4603} /* (24, 23, 8) {real, imag} */,
  {32'hc14afbc0, 32'h41aac09f} /* (24, 23, 7) {real, imag} */,
  {32'hc2d13736, 32'h4304b6c8} /* (24, 23, 6) {real, imag} */,
  {32'h4304d756, 32'h42c1fc15} /* (24, 23, 5) {real, imag} */,
  {32'hc326d0c5, 32'hc1ce6c5a} /* (24, 23, 4) {real, imag} */,
  {32'hc2bb865c, 32'hc19b8ca6} /* (24, 23, 3) {real, imag} */,
  {32'h44850fde, 32'h43418478} /* (24, 23, 2) {real, imag} */,
  {32'hc529e172, 32'hc3bbc3f2} /* (24, 23, 1) {real, imag} */,
  {32'hc529c570, 32'h00000000} /* (24, 23, 0) {real, imag} */,
  {32'hc50a861b, 32'h438405c5} /* (24, 22, 31) {real, imag} */,
  {32'h445cede4, 32'hc27331d8} /* (24, 22, 30) {real, imag} */,
  {32'hc0c0cc30, 32'h42894662} /* (24, 22, 29) {real, imag} */,
  {32'hc36fd172, 32'h43091f6b} /* (24, 22, 28) {real, imag} */,
  {32'h4389f72d, 32'hc2d9748a} /* (24, 22, 27) {real, imag} */,
  {32'hc303ea2a, 32'hc2c3df77} /* (24, 22, 26) {real, imag} */,
  {32'hc207b0f8, 32'h41f425aa} /* (24, 22, 25) {real, imag} */,
  {32'h41dd57d2, 32'hc1da7a41} /* (24, 22, 24) {real, imag} */,
  {32'hc15b5f50, 32'hc217fc99} /* (24, 22, 23) {real, imag} */,
  {32'hc20bf15e, 32'hc08954c4} /* (24, 22, 22) {real, imag} */,
  {32'hc2151428, 32'hc145ee96} /* (24, 22, 21) {real, imag} */,
  {32'h41c8e124, 32'h41dfc524} /* (24, 22, 20) {real, imag} */,
  {32'hc1dec561, 32'h42169040} /* (24, 22, 19) {real, imag} */,
  {32'h416acc5c, 32'h424c679c} /* (24, 22, 18) {real, imag} */,
  {32'h4288f0a1, 32'hc28a1499} /* (24, 22, 17) {real, imag} */,
  {32'hc1c364a4, 32'h00000000} /* (24, 22, 16) {real, imag} */,
  {32'h4288f0a1, 32'h428a1499} /* (24, 22, 15) {real, imag} */,
  {32'h416acc5c, 32'hc24c679c} /* (24, 22, 14) {real, imag} */,
  {32'hc1dec561, 32'hc2169040} /* (24, 22, 13) {real, imag} */,
  {32'h41c8e124, 32'hc1dfc524} /* (24, 22, 12) {real, imag} */,
  {32'hc2151428, 32'h4145ee96} /* (24, 22, 11) {real, imag} */,
  {32'hc20bf15e, 32'h408954c4} /* (24, 22, 10) {real, imag} */,
  {32'hc15b5f50, 32'h4217fc99} /* (24, 22, 9) {real, imag} */,
  {32'h41dd57d2, 32'h41da7a41} /* (24, 22, 8) {real, imag} */,
  {32'hc207b0f8, 32'hc1f425aa} /* (24, 22, 7) {real, imag} */,
  {32'hc303ea2a, 32'h42c3df77} /* (24, 22, 6) {real, imag} */,
  {32'h4389f72d, 32'h42d9748a} /* (24, 22, 5) {real, imag} */,
  {32'hc36fd172, 32'hc3091f6b} /* (24, 22, 4) {real, imag} */,
  {32'hc0c0cc30, 32'hc2894662} /* (24, 22, 3) {real, imag} */,
  {32'h445cede4, 32'h427331d8} /* (24, 22, 2) {real, imag} */,
  {32'hc50a861b, 32'hc38405c5} /* (24, 22, 1) {real, imag} */,
  {32'hc4f34d36, 32'h00000000} /* (24, 22, 0) {real, imag} */,
  {32'hc46602f0, 32'h42d62940} /* (24, 21, 31) {real, imag} */,
  {32'h43c5ebe7, 32'hc2d151ee} /* (24, 21, 30) {real, imag} */,
  {32'h422e1d4d, 32'h42badc45} /* (24, 21, 29) {real, imag} */,
  {32'h4237dce8, 32'h3fc9c200} /* (24, 21, 28) {real, imag} */,
  {32'h43261baa, 32'h4283890d} /* (24, 21, 27) {real, imag} */,
  {32'h4124fc9d, 32'h42e880a4} /* (24, 21, 26) {real, imag} */,
  {32'h42358709, 32'hc2a56231} /* (24, 21, 25) {real, imag} */,
  {32'hc1bc2b36, 32'h42219f17} /* (24, 21, 24) {real, imag} */,
  {32'hc31ca07c, 32'h41b14c08} /* (24, 21, 23) {real, imag} */,
  {32'h3fad8b68, 32'hc2813ebd} /* (24, 21, 22) {real, imag} */,
  {32'hc2fd67de, 32'h4154964f} /* (24, 21, 21) {real, imag} */,
  {32'h41ea8528, 32'h40933610} /* (24, 21, 20) {real, imag} */,
  {32'hc069d1e4, 32'hc12f6052} /* (24, 21, 19) {real, imag} */,
  {32'h422ed539, 32'h422fbe7c} /* (24, 21, 18) {real, imag} */,
  {32'hc1ad782e, 32'h411f1eec} /* (24, 21, 17) {real, imag} */,
  {32'h42216a5f, 32'h00000000} /* (24, 21, 16) {real, imag} */,
  {32'hc1ad782e, 32'hc11f1eec} /* (24, 21, 15) {real, imag} */,
  {32'h422ed539, 32'hc22fbe7c} /* (24, 21, 14) {real, imag} */,
  {32'hc069d1e4, 32'h412f6052} /* (24, 21, 13) {real, imag} */,
  {32'h41ea8528, 32'hc0933610} /* (24, 21, 12) {real, imag} */,
  {32'hc2fd67de, 32'hc154964f} /* (24, 21, 11) {real, imag} */,
  {32'h3fad8b68, 32'h42813ebd} /* (24, 21, 10) {real, imag} */,
  {32'hc31ca07c, 32'hc1b14c08} /* (24, 21, 9) {real, imag} */,
  {32'hc1bc2b36, 32'hc2219f17} /* (24, 21, 8) {real, imag} */,
  {32'h42358709, 32'h42a56231} /* (24, 21, 7) {real, imag} */,
  {32'h4124fc9d, 32'hc2e880a4} /* (24, 21, 6) {real, imag} */,
  {32'h43261baa, 32'hc283890d} /* (24, 21, 5) {real, imag} */,
  {32'h4237dce8, 32'hbfc9c200} /* (24, 21, 4) {real, imag} */,
  {32'h422e1d4d, 32'hc2badc45} /* (24, 21, 3) {real, imag} */,
  {32'h43c5ebe7, 32'h42d151ee} /* (24, 21, 2) {real, imag} */,
  {32'hc46602f0, 32'hc2d62940} /* (24, 21, 1) {real, imag} */,
  {32'hc4471abb, 32'h00000000} /* (24, 21, 0) {real, imag} */,
  {32'h44311f59, 32'hc3537cdc} /* (24, 20, 31) {real, imag} */,
  {32'hc3c8b2ec, 32'h42790f2c} /* (24, 20, 30) {real, imag} */,
  {32'h4298a550, 32'h43168d43} /* (24, 20, 29) {real, imag} */,
  {32'h4316e454, 32'hc312695d} /* (24, 20, 28) {real, imag} */,
  {32'hc2a02581, 32'h42b1cd76} /* (24, 20, 27) {real, imag} */,
  {32'h428bbc48, 32'h4227e60e} /* (24, 20, 26) {real, imag} */,
  {32'h42bf0696, 32'hc320b502} /* (24, 20, 25) {real, imag} */,
  {32'hc2dd47d9, 32'h424b33c6} /* (24, 20, 24) {real, imag} */,
  {32'hc2ab7ba0, 32'h430b400b} /* (24, 20, 23) {real, imag} */,
  {32'h42597ffc, 32'hc23bf132} /* (24, 20, 22) {real, imag} */,
  {32'h4269f585, 32'h42b0ae92} /* (24, 20, 21) {real, imag} */,
  {32'hc236782f, 32'hc220b746} /* (24, 20, 20) {real, imag} */,
  {32'hc2cf2f3e, 32'hc2a043f6} /* (24, 20, 19) {real, imag} */,
  {32'h428f0c92, 32'h418f2650} /* (24, 20, 18) {real, imag} */,
  {32'hc1cb7218, 32'h40d2e570} /* (24, 20, 17) {real, imag} */,
  {32'h41e3ad3e, 32'h00000000} /* (24, 20, 16) {real, imag} */,
  {32'hc1cb7218, 32'hc0d2e570} /* (24, 20, 15) {real, imag} */,
  {32'h428f0c92, 32'hc18f2650} /* (24, 20, 14) {real, imag} */,
  {32'hc2cf2f3e, 32'h42a043f6} /* (24, 20, 13) {real, imag} */,
  {32'hc236782f, 32'h4220b746} /* (24, 20, 12) {real, imag} */,
  {32'h4269f585, 32'hc2b0ae92} /* (24, 20, 11) {real, imag} */,
  {32'h42597ffc, 32'h423bf132} /* (24, 20, 10) {real, imag} */,
  {32'hc2ab7ba0, 32'hc30b400b} /* (24, 20, 9) {real, imag} */,
  {32'hc2dd47d9, 32'hc24b33c6} /* (24, 20, 8) {real, imag} */,
  {32'h42bf0696, 32'h4320b502} /* (24, 20, 7) {real, imag} */,
  {32'h428bbc48, 32'hc227e60e} /* (24, 20, 6) {real, imag} */,
  {32'hc2a02581, 32'hc2b1cd76} /* (24, 20, 5) {real, imag} */,
  {32'h4316e454, 32'h4312695d} /* (24, 20, 4) {real, imag} */,
  {32'h4298a550, 32'hc3168d43} /* (24, 20, 3) {real, imag} */,
  {32'hc3c8b2ec, 32'hc2790f2c} /* (24, 20, 2) {real, imag} */,
  {32'h44311f59, 32'h43537cdc} /* (24, 20, 1) {real, imag} */,
  {32'h43b768c6, 32'h00000000} /* (24, 20, 0) {real, imag} */,
  {32'h44c5b83a, 32'hc34443f8} /* (24, 19, 31) {real, imag} */,
  {32'hc44a3ac8, 32'h42ca1658} /* (24, 19, 30) {real, imag} */,
  {32'h4213ec54, 32'h42847107} /* (24, 19, 29) {real, imag} */,
  {32'h43436692, 32'hc3381637} /* (24, 19, 28) {real, imag} */,
  {32'hc30f7817, 32'h42f70c11} /* (24, 19, 27) {real, imag} */,
  {32'h42952ba0, 32'hc2165d93} /* (24, 19, 26) {real, imag} */,
  {32'h42541370, 32'h411d7637} /* (24, 19, 25) {real, imag} */,
  {32'hc334a3f4, 32'h42b94183} /* (24, 19, 24) {real, imag} */,
  {32'hc23fcb9b, 32'h3feb5310} /* (24, 19, 23) {real, imag} */,
  {32'h3f96b580, 32'h427f9728} /* (24, 19, 22) {real, imag} */,
  {32'h415e6653, 32'h4229ffdb} /* (24, 19, 21) {real, imag} */,
  {32'h418897c8, 32'hc1d50525} /* (24, 19, 20) {real, imag} */,
  {32'hc248dd06, 32'hc20ea6ea} /* (24, 19, 19) {real, imag} */,
  {32'hc20548aa, 32'h42371039} /* (24, 19, 18) {real, imag} */,
  {32'h42043c4c, 32'hc2595b1e} /* (24, 19, 17) {real, imag} */,
  {32'h40e9ef48, 32'h00000000} /* (24, 19, 16) {real, imag} */,
  {32'h42043c4c, 32'h42595b1e} /* (24, 19, 15) {real, imag} */,
  {32'hc20548aa, 32'hc2371039} /* (24, 19, 14) {real, imag} */,
  {32'hc248dd06, 32'h420ea6ea} /* (24, 19, 13) {real, imag} */,
  {32'h418897c8, 32'h41d50525} /* (24, 19, 12) {real, imag} */,
  {32'h415e6653, 32'hc229ffdb} /* (24, 19, 11) {real, imag} */,
  {32'h3f96b580, 32'hc27f9728} /* (24, 19, 10) {real, imag} */,
  {32'hc23fcb9b, 32'hbfeb5310} /* (24, 19, 9) {real, imag} */,
  {32'hc334a3f4, 32'hc2b94183} /* (24, 19, 8) {real, imag} */,
  {32'h42541370, 32'hc11d7637} /* (24, 19, 7) {real, imag} */,
  {32'h42952ba0, 32'h42165d93} /* (24, 19, 6) {real, imag} */,
  {32'hc30f7817, 32'hc2f70c11} /* (24, 19, 5) {real, imag} */,
  {32'h43436692, 32'h43381637} /* (24, 19, 4) {real, imag} */,
  {32'h4213ec54, 32'hc2847107} /* (24, 19, 3) {real, imag} */,
  {32'hc44a3ac8, 32'hc2ca1658} /* (24, 19, 2) {real, imag} */,
  {32'h44c5b83a, 32'h434443f8} /* (24, 19, 1) {real, imag} */,
  {32'h448972b3, 32'h00000000} /* (24, 19, 0) {real, imag} */,
  {32'h45084958, 32'hc37c266c} /* (24, 18, 31) {real, imag} */,
  {32'hc4514738, 32'h424d3806} /* (24, 18, 30) {real, imag} */,
  {32'h4315ccfe, 32'h40c8c1c0} /* (24, 18, 29) {real, imag} */,
  {32'h43778412, 32'hc354fc58} /* (24, 18, 28) {real, imag} */,
  {32'hc343802c, 32'h42a8c7dc} /* (24, 18, 27) {real, imag} */,
  {32'h42b88ff4, 32'hc282dc49} /* (24, 18, 26) {real, imag} */,
  {32'hc2916d1c, 32'h416c6e60} /* (24, 18, 25) {real, imag} */,
  {32'hc262e040, 32'h432838bc} /* (24, 18, 24) {real, imag} */,
  {32'h423cfc90, 32'hc1bdb7e8} /* (24, 18, 23) {real, imag} */,
  {32'h4251a4c6, 32'hc30aa28e} /* (24, 18, 22) {real, imag} */,
  {32'hc304c81d, 32'h43135481} /* (24, 18, 21) {real, imag} */,
  {32'h42a06a4a, 32'hc260ddd4} /* (24, 18, 20) {real, imag} */,
  {32'hc1ee9876, 32'h4200a9e4} /* (24, 18, 19) {real, imag} */,
  {32'h412fa871, 32'h428e3306} /* (24, 18, 18) {real, imag} */,
  {32'hc25d9e18, 32'hc146462f} /* (24, 18, 17) {real, imag} */,
  {32'hc1558a50, 32'h00000000} /* (24, 18, 16) {real, imag} */,
  {32'hc25d9e18, 32'h4146462f} /* (24, 18, 15) {real, imag} */,
  {32'h412fa871, 32'hc28e3306} /* (24, 18, 14) {real, imag} */,
  {32'hc1ee9876, 32'hc200a9e4} /* (24, 18, 13) {real, imag} */,
  {32'h42a06a4a, 32'h4260ddd4} /* (24, 18, 12) {real, imag} */,
  {32'hc304c81d, 32'hc3135481} /* (24, 18, 11) {real, imag} */,
  {32'h4251a4c6, 32'h430aa28e} /* (24, 18, 10) {real, imag} */,
  {32'h423cfc90, 32'h41bdb7e8} /* (24, 18, 9) {real, imag} */,
  {32'hc262e040, 32'hc32838bc} /* (24, 18, 8) {real, imag} */,
  {32'hc2916d1c, 32'hc16c6e60} /* (24, 18, 7) {real, imag} */,
  {32'h42b88ff4, 32'h4282dc49} /* (24, 18, 6) {real, imag} */,
  {32'hc343802c, 32'hc2a8c7dc} /* (24, 18, 5) {real, imag} */,
  {32'h43778412, 32'h4354fc58} /* (24, 18, 4) {real, imag} */,
  {32'h4315ccfe, 32'hc0c8c1c0} /* (24, 18, 3) {real, imag} */,
  {32'hc4514738, 32'hc24d3806} /* (24, 18, 2) {real, imag} */,
  {32'h45084958, 32'h437c266c} /* (24, 18, 1) {real, imag} */,
  {32'h44cb0dd9, 32'h00000000} /* (24, 18, 0) {real, imag} */,
  {32'h45286346, 32'hc3ba94a6} /* (24, 17, 31) {real, imag} */,
  {32'hc4576bb6, 32'h434d8d3d} /* (24, 17, 30) {real, imag} */,
  {32'h42b2093e, 32'h423a8210} /* (24, 17, 29) {real, imag} */,
  {32'h43716fce, 32'hc2d031b2} /* (24, 17, 28) {real, imag} */,
  {32'hc2e32c00, 32'h4201fd6e} /* (24, 17, 27) {real, imag} */,
  {32'h4298fa0a, 32'h425bea1c} /* (24, 17, 26) {real, imag} */,
  {32'h42a29936, 32'hc08abce4} /* (24, 17, 25) {real, imag} */,
  {32'h4224e1a6, 32'h41c2604c} /* (24, 17, 24) {real, imag} */,
  {32'h40ad7e2c, 32'hc203c173} /* (24, 17, 23) {real, imag} */,
  {32'h41dd90a8, 32'h40b1270c} /* (24, 17, 22) {real, imag} */,
  {32'h41e0dc80, 32'h42f6a1b5} /* (24, 17, 21) {real, imag} */,
  {32'h41889737, 32'h41e0bf06} /* (24, 17, 20) {real, imag} */,
  {32'hc084539c, 32'h421ab4cd} /* (24, 17, 19) {real, imag} */,
  {32'h42be4488, 32'hc18b63d0} /* (24, 17, 18) {real, imag} */,
  {32'hc17aded4, 32'hc13b5bbe} /* (24, 17, 17) {real, imag} */,
  {32'hc1f14771, 32'h00000000} /* (24, 17, 16) {real, imag} */,
  {32'hc17aded4, 32'h413b5bbe} /* (24, 17, 15) {real, imag} */,
  {32'h42be4488, 32'h418b63d0} /* (24, 17, 14) {real, imag} */,
  {32'hc084539c, 32'hc21ab4cd} /* (24, 17, 13) {real, imag} */,
  {32'h41889737, 32'hc1e0bf06} /* (24, 17, 12) {real, imag} */,
  {32'h41e0dc80, 32'hc2f6a1b5} /* (24, 17, 11) {real, imag} */,
  {32'h41dd90a8, 32'hc0b1270c} /* (24, 17, 10) {real, imag} */,
  {32'h40ad7e2c, 32'h4203c173} /* (24, 17, 9) {real, imag} */,
  {32'h4224e1a6, 32'hc1c2604c} /* (24, 17, 8) {real, imag} */,
  {32'h42a29936, 32'h408abce4} /* (24, 17, 7) {real, imag} */,
  {32'h4298fa0a, 32'hc25bea1c} /* (24, 17, 6) {real, imag} */,
  {32'hc2e32c00, 32'hc201fd6e} /* (24, 17, 5) {real, imag} */,
  {32'h43716fce, 32'h42d031b2} /* (24, 17, 4) {real, imag} */,
  {32'h42b2093e, 32'hc23a8210} /* (24, 17, 3) {real, imag} */,
  {32'hc4576bb6, 32'hc34d8d3d} /* (24, 17, 2) {real, imag} */,
  {32'h45286346, 32'h43ba94a6} /* (24, 17, 1) {real, imag} */,
  {32'h44e402eb, 32'h00000000} /* (24, 17, 0) {real, imag} */,
  {32'h45389e85, 32'hc36b8300} /* (24, 16, 31) {real, imag} */,
  {32'hc468f100, 32'h43b2bd8a} /* (24, 16, 30) {real, imag} */,
  {32'hc18323f8, 32'h424b1b94} /* (24, 16, 29) {real, imag} */,
  {32'h43a77233, 32'hc33ce9a2} /* (24, 16, 28) {real, imag} */,
  {32'hc385d903, 32'hc1e33589} /* (24, 16, 27) {real, imag} */,
  {32'h4227c0e8, 32'h422d9848} /* (24, 16, 26) {real, imag} */,
  {32'h42b00872, 32'hc0cf771c} /* (24, 16, 25) {real, imag} */,
  {32'hc2e8cd90, 32'h42d26a5d} /* (24, 16, 24) {real, imag} */,
  {32'h427b71d3, 32'hbb87d800} /* (24, 16, 23) {real, imag} */,
  {32'hc29ac810, 32'h4254c88d} /* (24, 16, 22) {real, imag} */,
  {32'hc1938fc6, 32'h42d59cae} /* (24, 16, 21) {real, imag} */,
  {32'h40e1b30b, 32'hc1f48737} /* (24, 16, 20) {real, imag} */,
  {32'h41995e28, 32'hc19e2a2e} /* (24, 16, 19) {real, imag} */,
  {32'h41bbcf1a, 32'hc142011b} /* (24, 16, 18) {real, imag} */,
  {32'h4226b8a3, 32'h424e5148} /* (24, 16, 17) {real, imag} */,
  {32'hc20d51b8, 32'h00000000} /* (24, 16, 16) {real, imag} */,
  {32'h4226b8a3, 32'hc24e5148} /* (24, 16, 15) {real, imag} */,
  {32'h41bbcf1a, 32'h4142011b} /* (24, 16, 14) {real, imag} */,
  {32'h41995e28, 32'h419e2a2e} /* (24, 16, 13) {real, imag} */,
  {32'h40e1b30b, 32'h41f48737} /* (24, 16, 12) {real, imag} */,
  {32'hc1938fc6, 32'hc2d59cae} /* (24, 16, 11) {real, imag} */,
  {32'hc29ac810, 32'hc254c88d} /* (24, 16, 10) {real, imag} */,
  {32'h427b71d3, 32'h3b87d800} /* (24, 16, 9) {real, imag} */,
  {32'hc2e8cd90, 32'hc2d26a5d} /* (24, 16, 8) {real, imag} */,
  {32'h42b00872, 32'h40cf771c} /* (24, 16, 7) {real, imag} */,
  {32'h4227c0e8, 32'hc22d9848} /* (24, 16, 6) {real, imag} */,
  {32'hc385d903, 32'h41e33589} /* (24, 16, 5) {real, imag} */,
  {32'h43a77233, 32'h433ce9a2} /* (24, 16, 4) {real, imag} */,
  {32'hc18323f8, 32'hc24b1b94} /* (24, 16, 3) {real, imag} */,
  {32'hc468f100, 32'hc3b2bd8a} /* (24, 16, 2) {real, imag} */,
  {32'h45389e85, 32'h436b8300} /* (24, 16, 1) {real, imag} */,
  {32'h44f7c388, 32'h00000000} /* (24, 16, 0) {real, imag} */,
  {32'h453350f2, 32'hc32f4e15} /* (24, 15, 31) {real, imag} */,
  {32'hc465b0ca, 32'h438776fe} /* (24, 15, 30) {real, imag} */,
  {32'hc26cc200, 32'h40e2cf40} /* (24, 15, 29) {real, imag} */,
  {32'h43311eca, 32'hc260824c} /* (24, 15, 28) {real, imag} */,
  {32'hc35db7f2, 32'h41d1e001} /* (24, 15, 27) {real, imag} */,
  {32'hc0ba61f8, 32'h428d7187} /* (24, 15, 26) {real, imag} */,
  {32'h41346ddc, 32'hbf97c870} /* (24, 15, 25) {real, imag} */,
  {32'hc2b27213, 32'h410540c1} /* (24, 15, 24) {real, imag} */,
  {32'hc04aa878, 32'hc286716a} /* (24, 15, 23) {real, imag} */,
  {32'hc1994240, 32'h418c96e5} /* (24, 15, 22) {real, imag} */,
  {32'h41f89af0, 32'h42108b5a} /* (24, 15, 21) {real, imag} */,
  {32'hc16fcdda, 32'hc2945a88} /* (24, 15, 20) {real, imag} */,
  {32'h423edc34, 32'h42e3a962} /* (24, 15, 19) {real, imag} */,
  {32'h400035e0, 32'h4132447b} /* (24, 15, 18) {real, imag} */,
  {32'h4197887a, 32'h4125e40e} /* (24, 15, 17) {real, imag} */,
  {32'hc1e7f9f3, 32'h00000000} /* (24, 15, 16) {real, imag} */,
  {32'h4197887a, 32'hc125e40e} /* (24, 15, 15) {real, imag} */,
  {32'h400035e0, 32'hc132447b} /* (24, 15, 14) {real, imag} */,
  {32'h423edc34, 32'hc2e3a962} /* (24, 15, 13) {real, imag} */,
  {32'hc16fcdda, 32'h42945a88} /* (24, 15, 12) {real, imag} */,
  {32'h41f89af0, 32'hc2108b5a} /* (24, 15, 11) {real, imag} */,
  {32'hc1994240, 32'hc18c96e5} /* (24, 15, 10) {real, imag} */,
  {32'hc04aa878, 32'h4286716a} /* (24, 15, 9) {real, imag} */,
  {32'hc2b27213, 32'hc10540c1} /* (24, 15, 8) {real, imag} */,
  {32'h41346ddc, 32'h3f97c870} /* (24, 15, 7) {real, imag} */,
  {32'hc0ba61f8, 32'hc28d7187} /* (24, 15, 6) {real, imag} */,
  {32'hc35db7f2, 32'hc1d1e001} /* (24, 15, 5) {real, imag} */,
  {32'h43311eca, 32'h4260824c} /* (24, 15, 4) {real, imag} */,
  {32'hc26cc200, 32'hc0e2cf40} /* (24, 15, 3) {real, imag} */,
  {32'hc465b0ca, 32'hc38776fe} /* (24, 15, 2) {real, imag} */,
  {32'h453350f2, 32'h432f4e15} /* (24, 15, 1) {real, imag} */,
  {32'h44ede86d, 32'h00000000} /* (24, 15, 0) {real, imag} */,
  {32'h452b539c, 32'hc2f0d248} /* (24, 14, 31) {real, imag} */,
  {32'hc48ffb0f, 32'h4383294c} /* (24, 14, 30) {real, imag} */,
  {32'hc22b835a, 32'h42cd469e} /* (24, 14, 29) {real, imag} */,
  {32'h4325c904, 32'hc33b8e86} /* (24, 14, 28) {real, imag} */,
  {32'hc3367528, 32'h4240efc0} /* (24, 14, 27) {real, imag} */,
  {32'hc11b06a4, 32'h3fdf43f0} /* (24, 14, 26) {real, imag} */,
  {32'h431049e4, 32'hc28b63a8} /* (24, 14, 25) {real, imag} */,
  {32'hc1e13b08, 32'hc17fc818} /* (24, 14, 24) {real, imag} */,
  {32'hc1c3528f, 32'h4286a725} /* (24, 14, 23) {real, imag} */,
  {32'hc22614c6, 32'h3f066800} /* (24, 14, 22) {real, imag} */,
  {32'h425a7ba3, 32'hc1fa3a08} /* (24, 14, 21) {real, imag} */,
  {32'hc25e6298, 32'hc249aade} /* (24, 14, 20) {real, imag} */,
  {32'hc0d1d1b8, 32'h424ec6f6} /* (24, 14, 19) {real, imag} */,
  {32'h41548331, 32'h40ca9028} /* (24, 14, 18) {real, imag} */,
  {32'hc1bd1ce9, 32'hc098adee} /* (24, 14, 17) {real, imag} */,
  {32'h426cd196, 32'h00000000} /* (24, 14, 16) {real, imag} */,
  {32'hc1bd1ce9, 32'h4098adee} /* (24, 14, 15) {real, imag} */,
  {32'h41548331, 32'hc0ca9028} /* (24, 14, 14) {real, imag} */,
  {32'hc0d1d1b8, 32'hc24ec6f6} /* (24, 14, 13) {real, imag} */,
  {32'hc25e6298, 32'h4249aade} /* (24, 14, 12) {real, imag} */,
  {32'h425a7ba3, 32'h41fa3a08} /* (24, 14, 11) {real, imag} */,
  {32'hc22614c6, 32'hbf066800} /* (24, 14, 10) {real, imag} */,
  {32'hc1c3528f, 32'hc286a725} /* (24, 14, 9) {real, imag} */,
  {32'hc1e13b08, 32'h417fc818} /* (24, 14, 8) {real, imag} */,
  {32'h431049e4, 32'h428b63a8} /* (24, 14, 7) {real, imag} */,
  {32'hc11b06a4, 32'hbfdf43f0} /* (24, 14, 6) {real, imag} */,
  {32'hc3367528, 32'hc240efc0} /* (24, 14, 5) {real, imag} */,
  {32'h4325c904, 32'h433b8e86} /* (24, 14, 4) {real, imag} */,
  {32'hc22b835a, 32'hc2cd469e} /* (24, 14, 3) {real, imag} */,
  {32'hc48ffb0f, 32'hc383294c} /* (24, 14, 2) {real, imag} */,
  {32'h452b539c, 32'h42f0d248} /* (24, 14, 1) {real, imag} */,
  {32'h44ef6213, 32'h00000000} /* (24, 14, 0) {real, imag} */,
  {32'h451829df, 32'h406ea200} /* (24, 13, 31) {real, imag} */,
  {32'hc48e5552, 32'h432e2050} /* (24, 13, 30) {real, imag} */,
  {32'hc32b7ed3, 32'h42523cbe} /* (24, 13, 29) {real, imag} */,
  {32'h431db460, 32'hc379cf2b} /* (24, 13, 28) {real, imag} */,
  {32'hc36eac33, 32'h42587a6a} /* (24, 13, 27) {real, imag} */,
  {32'h42480351, 32'h40aeefe8} /* (24, 13, 26) {real, imag} */,
  {32'h42f0eaf8, 32'hc170e155} /* (24, 13, 25) {real, imag} */,
  {32'h42cae87b, 32'h3ffc01c0} /* (24, 13, 24) {real, imag} */,
  {32'hc2b3667a, 32'hc2578ee4} /* (24, 13, 23) {real, imag} */,
  {32'hc1159908, 32'h424969ca} /* (24, 13, 22) {real, imag} */,
  {32'h4184385a, 32'hc14dc259} /* (24, 13, 21) {real, imag} */,
  {32'hc0e48ec0, 32'hc27e5bbe} /* (24, 13, 20) {real, imag} */,
  {32'hc0a7f430, 32'h41fb87cc} /* (24, 13, 19) {real, imag} */,
  {32'h40423038, 32'h42d9e124} /* (24, 13, 18) {real, imag} */,
  {32'hc13da112, 32'hc1bbfae0} /* (24, 13, 17) {real, imag} */,
  {32'hc1808992, 32'h00000000} /* (24, 13, 16) {real, imag} */,
  {32'hc13da112, 32'h41bbfae0} /* (24, 13, 15) {real, imag} */,
  {32'h40423038, 32'hc2d9e124} /* (24, 13, 14) {real, imag} */,
  {32'hc0a7f430, 32'hc1fb87cc} /* (24, 13, 13) {real, imag} */,
  {32'hc0e48ec0, 32'h427e5bbe} /* (24, 13, 12) {real, imag} */,
  {32'h4184385a, 32'h414dc259} /* (24, 13, 11) {real, imag} */,
  {32'hc1159908, 32'hc24969ca} /* (24, 13, 10) {real, imag} */,
  {32'hc2b3667a, 32'h42578ee4} /* (24, 13, 9) {real, imag} */,
  {32'h42cae87b, 32'hbffc01c0} /* (24, 13, 8) {real, imag} */,
  {32'h42f0eaf8, 32'h4170e155} /* (24, 13, 7) {real, imag} */,
  {32'h42480351, 32'hc0aeefe8} /* (24, 13, 6) {real, imag} */,
  {32'hc36eac33, 32'hc2587a6a} /* (24, 13, 5) {real, imag} */,
  {32'h431db460, 32'h4379cf2b} /* (24, 13, 4) {real, imag} */,
  {32'hc32b7ed3, 32'hc2523cbe} /* (24, 13, 3) {real, imag} */,
  {32'hc48e5552, 32'hc32e2050} /* (24, 13, 2) {real, imag} */,
  {32'h451829df, 32'hc06ea200} /* (24, 13, 1) {real, imag} */,
  {32'h44d69d05, 32'h00000000} /* (24, 13, 0) {real, imag} */,
  {32'h44f8daea, 32'h43580884} /* (24, 12, 31) {real, imag} */,
  {32'hc483e80d, 32'hc1228a70} /* (24, 12, 30) {real, imag} */,
  {32'hc238ac65, 32'h42b79bbc} /* (24, 12, 29) {real, imag} */,
  {32'h433f00c0, 32'hc2c159c6} /* (24, 12, 28) {real, imag} */,
  {32'hc2d14cd7, 32'h4336f08b} /* (24, 12, 27) {real, imag} */,
  {32'h41993c3a, 32'hc243bbd0} /* (24, 12, 26) {real, imag} */,
  {32'h42dbc6d6, 32'h420c69ad} /* (24, 12, 25) {real, imag} */,
  {32'hbfa31700, 32'h42ccd9f5} /* (24, 12, 24) {real, imag} */,
  {32'hc2825024, 32'hc2d3b99a} /* (24, 12, 23) {real, imag} */,
  {32'hc01530e8, 32'h42aecf3b} /* (24, 12, 22) {real, imag} */,
  {32'hc0c2a158, 32'h419d4822} /* (24, 12, 21) {real, imag} */,
  {32'h4268cf65, 32'h420ac2f2} /* (24, 12, 20) {real, imag} */,
  {32'h41cc7a48, 32'h429af994} /* (24, 12, 19) {real, imag} */,
  {32'hc2442b76, 32'h42e2d434} /* (24, 12, 18) {real, imag} */,
  {32'hc28e52de, 32'hc2b25341} /* (24, 12, 17) {real, imag} */,
  {32'h42c6112e, 32'h00000000} /* (24, 12, 16) {real, imag} */,
  {32'hc28e52de, 32'h42b25341} /* (24, 12, 15) {real, imag} */,
  {32'hc2442b76, 32'hc2e2d434} /* (24, 12, 14) {real, imag} */,
  {32'h41cc7a48, 32'hc29af994} /* (24, 12, 13) {real, imag} */,
  {32'h4268cf65, 32'hc20ac2f2} /* (24, 12, 12) {real, imag} */,
  {32'hc0c2a158, 32'hc19d4822} /* (24, 12, 11) {real, imag} */,
  {32'hc01530e8, 32'hc2aecf3b} /* (24, 12, 10) {real, imag} */,
  {32'hc2825024, 32'h42d3b99a} /* (24, 12, 9) {real, imag} */,
  {32'hbfa31700, 32'hc2ccd9f5} /* (24, 12, 8) {real, imag} */,
  {32'h42dbc6d6, 32'hc20c69ad} /* (24, 12, 7) {real, imag} */,
  {32'h41993c3a, 32'h4243bbd0} /* (24, 12, 6) {real, imag} */,
  {32'hc2d14cd7, 32'hc336f08b} /* (24, 12, 5) {real, imag} */,
  {32'h433f00c0, 32'h42c159c6} /* (24, 12, 4) {real, imag} */,
  {32'hc238ac65, 32'hc2b79bbc} /* (24, 12, 3) {real, imag} */,
  {32'hc483e80d, 32'h41228a70} /* (24, 12, 2) {real, imag} */,
  {32'h44f8daea, 32'hc3580884} /* (24, 12, 1) {real, imag} */,
  {32'h4491b764, 32'h00000000} /* (24, 12, 0) {real, imag} */,
  {32'h44737814, 32'h43afe7f0} /* (24, 11, 31) {real, imag} */,
  {32'hc44caa70, 32'hc24a9644} /* (24, 11, 30) {real, imag} */,
  {32'hc21fe157, 32'h4295eaab} /* (24, 11, 29) {real, imag} */,
  {32'h439dc889, 32'hc3698aec} /* (24, 11, 28) {real, imag} */,
  {32'h401a3d60, 32'h4225620e} /* (24, 11, 27) {real, imag} */,
  {32'hc0e6c92a, 32'h42bf33d4} /* (24, 11, 26) {real, imag} */,
  {32'hc2742053, 32'hc2809547} /* (24, 11, 25) {real, imag} */,
  {32'hc3164b53, 32'h4123c733} /* (24, 11, 24) {real, imag} */,
  {32'hc2a59b85, 32'h41d1af34} /* (24, 11, 23) {real, imag} */,
  {32'h41fc0c84, 32'hc11d2a86} /* (24, 11, 22) {real, imag} */,
  {32'hc15672e0, 32'h41ccd2d0} /* (24, 11, 21) {real, imag} */,
  {32'h41a26636, 32'h42c90a4a} /* (24, 11, 20) {real, imag} */,
  {32'hc2063211, 32'hc1dc5dcb} /* (24, 11, 19) {real, imag} */,
  {32'h429854f8, 32'hc0568c68} /* (24, 11, 18) {real, imag} */,
  {32'h41592489, 32'h42b31826} /* (24, 11, 17) {real, imag} */,
  {32'h42d2aadc, 32'h00000000} /* (24, 11, 16) {real, imag} */,
  {32'h41592489, 32'hc2b31826} /* (24, 11, 15) {real, imag} */,
  {32'h429854f8, 32'h40568c68} /* (24, 11, 14) {real, imag} */,
  {32'hc2063211, 32'h41dc5dcb} /* (24, 11, 13) {real, imag} */,
  {32'h41a26636, 32'hc2c90a4a} /* (24, 11, 12) {real, imag} */,
  {32'hc15672e0, 32'hc1ccd2d0} /* (24, 11, 11) {real, imag} */,
  {32'h41fc0c84, 32'h411d2a86} /* (24, 11, 10) {real, imag} */,
  {32'hc2a59b85, 32'hc1d1af34} /* (24, 11, 9) {real, imag} */,
  {32'hc3164b53, 32'hc123c733} /* (24, 11, 8) {real, imag} */,
  {32'hc2742053, 32'h42809547} /* (24, 11, 7) {real, imag} */,
  {32'hc0e6c92a, 32'hc2bf33d4} /* (24, 11, 6) {real, imag} */,
  {32'h401a3d60, 32'hc225620e} /* (24, 11, 5) {real, imag} */,
  {32'h439dc889, 32'h43698aec} /* (24, 11, 4) {real, imag} */,
  {32'hc21fe157, 32'hc295eaab} /* (24, 11, 3) {real, imag} */,
  {32'hc44caa70, 32'h424a9644} /* (24, 11, 2) {real, imag} */,
  {32'h44737814, 32'hc3afe7f0} /* (24, 11, 1) {real, imag} */,
  {32'h4412fe9f, 32'h00000000} /* (24, 11, 0) {real, imag} */,
  {32'hc420177b, 32'h441a0276} /* (24, 10, 31) {real, imag} */,
  {32'h40118a80, 32'hc32c4fe0} /* (24, 10, 30) {real, imag} */,
  {32'hc30aefaa, 32'h41636344} /* (24, 10, 29) {real, imag} */,
  {32'h42e5405c, 32'hc2f6b5aa} /* (24, 10, 28) {real, imag} */,
  {32'h42dca0d3, 32'hc20645fc} /* (24, 10, 27) {real, imag} */,
  {32'h423a0403, 32'h41c34ff4} /* (24, 10, 26) {real, imag} */,
  {32'h41fafd5f, 32'h42fa5e26} /* (24, 10, 25) {real, imag} */,
  {32'h419b721e, 32'hc1d186a5} /* (24, 10, 24) {real, imag} */,
  {32'hc29ff736, 32'h4201595f} /* (24, 10, 23) {real, imag} */,
  {32'hc1d61b65, 32'hc1b04525} /* (24, 10, 22) {real, imag} */,
  {32'hc22fe0e4, 32'hc297c74f} /* (24, 10, 21) {real, imag} */,
  {32'hc2b82a04, 32'hc2bc3c9f} /* (24, 10, 20) {real, imag} */,
  {32'h41ed3bd1, 32'hc301e6fc} /* (24, 10, 19) {real, imag} */,
  {32'hc11a3e00, 32'hc203afe8} /* (24, 10, 18) {real, imag} */,
  {32'hc1282b4a, 32'h4115f546} /* (24, 10, 17) {real, imag} */,
  {32'hc27c5456, 32'h00000000} /* (24, 10, 16) {real, imag} */,
  {32'hc1282b4a, 32'hc115f546} /* (24, 10, 15) {real, imag} */,
  {32'hc11a3e00, 32'h4203afe8} /* (24, 10, 14) {real, imag} */,
  {32'h41ed3bd1, 32'h4301e6fc} /* (24, 10, 13) {real, imag} */,
  {32'hc2b82a04, 32'h42bc3c9f} /* (24, 10, 12) {real, imag} */,
  {32'hc22fe0e4, 32'h4297c74f} /* (24, 10, 11) {real, imag} */,
  {32'hc1d61b65, 32'h41b04525} /* (24, 10, 10) {real, imag} */,
  {32'hc29ff736, 32'hc201595f} /* (24, 10, 9) {real, imag} */,
  {32'h419b721e, 32'h41d186a5} /* (24, 10, 8) {real, imag} */,
  {32'h41fafd5f, 32'hc2fa5e26} /* (24, 10, 7) {real, imag} */,
  {32'h423a0403, 32'hc1c34ff4} /* (24, 10, 6) {real, imag} */,
  {32'h42dca0d3, 32'h420645fc} /* (24, 10, 5) {real, imag} */,
  {32'h42e5405c, 32'h42f6b5aa} /* (24, 10, 4) {real, imag} */,
  {32'hc30aefaa, 32'hc1636344} /* (24, 10, 3) {real, imag} */,
  {32'h40118a80, 32'h432c4fe0} /* (24, 10, 2) {real, imag} */,
  {32'hc420177b, 32'hc41a0276} /* (24, 10, 1) {real, imag} */,
  {32'hc42c5009, 32'h00000000} /* (24, 10, 0) {real, imag} */,
  {32'hc4da16e0, 32'h446db447} /* (24, 9, 31) {real, imag} */,
  {32'h43fa7478, 32'hc3664fb0} /* (24, 9, 30) {real, imag} */,
  {32'hc04fd310, 32'hc1545974} /* (24, 9, 29) {real, imag} */,
  {32'hc2096680, 32'hc2a8f86c} /* (24, 9, 28) {real, imag} */,
  {32'h42c48646, 32'hc2c9259b} /* (24, 9, 27) {real, imag} */,
  {32'h4269a4e3, 32'hc13dba00} /* (24, 9, 26) {real, imag} */,
  {32'h41a28680, 32'h418dc55f} /* (24, 9, 25) {real, imag} */,
  {32'h4243753c, 32'h420b3c6e} /* (24, 9, 24) {real, imag} */,
  {32'h42959758, 32'h429a5656} /* (24, 9, 23) {real, imag} */,
  {32'h420e4db9, 32'hc1c55b13} /* (24, 9, 22) {real, imag} */,
  {32'hc2d927e0, 32'hc28afc1a} /* (24, 9, 21) {real, imag} */,
  {32'hc23e5ae1, 32'h421f27ac} /* (24, 9, 20) {real, imag} */,
  {32'h41d62d26, 32'hc2a06cf2} /* (24, 9, 19) {real, imag} */,
  {32'h42b5f3ed, 32'h3ee0b820} /* (24, 9, 18) {real, imag} */,
  {32'hc1910b40, 32'hc1dd3b35} /* (24, 9, 17) {real, imag} */,
  {32'h425f535b, 32'h00000000} /* (24, 9, 16) {real, imag} */,
  {32'hc1910b40, 32'h41dd3b35} /* (24, 9, 15) {real, imag} */,
  {32'h42b5f3ed, 32'hbee0b820} /* (24, 9, 14) {real, imag} */,
  {32'h41d62d26, 32'h42a06cf2} /* (24, 9, 13) {real, imag} */,
  {32'hc23e5ae1, 32'hc21f27ac} /* (24, 9, 12) {real, imag} */,
  {32'hc2d927e0, 32'h428afc1a} /* (24, 9, 11) {real, imag} */,
  {32'h420e4db9, 32'h41c55b13} /* (24, 9, 10) {real, imag} */,
  {32'h42959758, 32'hc29a5656} /* (24, 9, 9) {real, imag} */,
  {32'h4243753c, 32'hc20b3c6e} /* (24, 9, 8) {real, imag} */,
  {32'h41a28680, 32'hc18dc55f} /* (24, 9, 7) {real, imag} */,
  {32'h4269a4e3, 32'h413dba00} /* (24, 9, 6) {real, imag} */,
  {32'h42c48646, 32'h42c9259b} /* (24, 9, 5) {real, imag} */,
  {32'hc2096680, 32'h42a8f86c} /* (24, 9, 4) {real, imag} */,
  {32'hc04fd310, 32'h41545974} /* (24, 9, 3) {real, imag} */,
  {32'h43fa7478, 32'h43664fb0} /* (24, 9, 2) {real, imag} */,
  {32'hc4da16e0, 32'hc46db447} /* (24, 9, 1) {real, imag} */,
  {32'hc4e9481b, 32'h00000000} /* (24, 9, 0) {real, imag} */,
  {32'hc5120b28, 32'h4494d9d1} /* (24, 8, 31) {real, imag} */,
  {32'h44358c36, 32'hc3b9d678} /* (24, 8, 30) {real, imag} */,
  {32'h43057e3d, 32'h42b31102} /* (24, 8, 29) {real, imag} */,
  {32'hc3172f33, 32'h422293fd} /* (24, 8, 28) {real, imag} */,
  {32'h414930e8, 32'hc3401e0b} /* (24, 8, 27) {real, imag} */,
  {32'h429d4416, 32'hc309385a} /* (24, 8, 26) {real, imag} */,
  {32'h427bb1c4, 32'hc2e3f329} /* (24, 8, 25) {real, imag} */,
  {32'h42ec11df, 32'hc2413328} /* (24, 8, 24) {real, imag} */,
  {32'hc2cc06ff, 32'h41f6c6a2} /* (24, 8, 23) {real, imag} */,
  {32'h41c62402, 32'h41011420} /* (24, 8, 22) {real, imag} */,
  {32'h428af28d, 32'h425d1ac0} /* (24, 8, 21) {real, imag} */,
  {32'h42699ed9, 32'h41d14e1a} /* (24, 8, 20) {real, imag} */,
  {32'h4150f1d9, 32'h428fc793} /* (24, 8, 19) {real, imag} */,
  {32'h4263903c, 32'h411ccfe8} /* (24, 8, 18) {real, imag} */,
  {32'h424e1ea9, 32'h4240c937} /* (24, 8, 17) {real, imag} */,
  {32'h40c1ffb0, 32'h00000000} /* (24, 8, 16) {real, imag} */,
  {32'h424e1ea9, 32'hc240c937} /* (24, 8, 15) {real, imag} */,
  {32'h4263903c, 32'hc11ccfe8} /* (24, 8, 14) {real, imag} */,
  {32'h4150f1d9, 32'hc28fc793} /* (24, 8, 13) {real, imag} */,
  {32'h42699ed9, 32'hc1d14e1a} /* (24, 8, 12) {real, imag} */,
  {32'h428af28d, 32'hc25d1ac0} /* (24, 8, 11) {real, imag} */,
  {32'h41c62402, 32'hc1011420} /* (24, 8, 10) {real, imag} */,
  {32'hc2cc06ff, 32'hc1f6c6a2} /* (24, 8, 9) {real, imag} */,
  {32'h42ec11df, 32'h42413328} /* (24, 8, 8) {real, imag} */,
  {32'h427bb1c4, 32'h42e3f329} /* (24, 8, 7) {real, imag} */,
  {32'h429d4416, 32'h4309385a} /* (24, 8, 6) {real, imag} */,
  {32'h414930e8, 32'h43401e0b} /* (24, 8, 5) {real, imag} */,
  {32'hc3172f33, 32'hc22293fd} /* (24, 8, 4) {real, imag} */,
  {32'h43057e3d, 32'hc2b31102} /* (24, 8, 3) {real, imag} */,
  {32'h44358c36, 32'h43b9d678} /* (24, 8, 2) {real, imag} */,
  {32'hc5120b28, 32'hc494d9d1} /* (24, 8, 1) {real, imag} */,
  {32'hc521628e, 32'h00000000} /* (24, 8, 0) {real, imag} */,
  {32'hc525ab9f, 32'h44b5c158} /* (24, 7, 31) {real, imag} */,
  {32'h4427217a, 32'hc39e61da} /* (24, 7, 30) {real, imag} */,
  {32'h42d9cb72, 32'hc1e7881b} /* (24, 7, 29) {real, imag} */,
  {32'hc363e172, 32'h41a9675f} /* (24, 7, 28) {real, imag} */,
  {32'h432783c2, 32'hc20f7239} /* (24, 7, 27) {real, imag} */,
  {32'h42aaa0a8, 32'hc248f723} /* (24, 7, 26) {real, imag} */,
  {32'hc303b5e0, 32'hc18b736e} /* (24, 7, 25) {real, imag} */,
  {32'h42db72c5, 32'hc25ee4e6} /* (24, 7, 24) {real, imag} */,
  {32'hc2301335, 32'hc241aa24} /* (24, 7, 23) {real, imag} */,
  {32'h42cc6190, 32'h42a2e487} /* (24, 7, 22) {real, imag} */,
  {32'h41383a18, 32'hc2b0168f} /* (24, 7, 21) {real, imag} */,
  {32'hc2e2ad8a, 32'hc24480e8} /* (24, 7, 20) {real, imag} */,
  {32'h42286b2c, 32'hc1376a54} /* (24, 7, 19) {real, imag} */,
  {32'h401d7f90, 32'hc1e69474} /* (24, 7, 18) {real, imag} */,
  {32'hc1d378e9, 32'hc141af1d} /* (24, 7, 17) {real, imag} */,
  {32'h4096d75c, 32'h00000000} /* (24, 7, 16) {real, imag} */,
  {32'hc1d378e9, 32'h4141af1d} /* (24, 7, 15) {real, imag} */,
  {32'h401d7f90, 32'h41e69474} /* (24, 7, 14) {real, imag} */,
  {32'h42286b2c, 32'h41376a54} /* (24, 7, 13) {real, imag} */,
  {32'hc2e2ad8a, 32'h424480e8} /* (24, 7, 12) {real, imag} */,
  {32'h41383a18, 32'h42b0168f} /* (24, 7, 11) {real, imag} */,
  {32'h42cc6190, 32'hc2a2e487} /* (24, 7, 10) {real, imag} */,
  {32'hc2301335, 32'h4241aa24} /* (24, 7, 9) {real, imag} */,
  {32'h42db72c5, 32'h425ee4e6} /* (24, 7, 8) {real, imag} */,
  {32'hc303b5e0, 32'h418b736e} /* (24, 7, 7) {real, imag} */,
  {32'h42aaa0a8, 32'h4248f723} /* (24, 7, 6) {real, imag} */,
  {32'h432783c2, 32'h420f7239} /* (24, 7, 5) {real, imag} */,
  {32'hc363e172, 32'hc1a9675f} /* (24, 7, 4) {real, imag} */,
  {32'h42d9cb72, 32'h41e7881b} /* (24, 7, 3) {real, imag} */,
  {32'h4427217a, 32'h439e61da} /* (24, 7, 2) {real, imag} */,
  {32'hc525ab9f, 32'hc4b5c158} /* (24, 7, 1) {real, imag} */,
  {32'hc5483cf8, 32'h00000000} /* (24, 7, 0) {real, imag} */,
  {32'hc52d7c4b, 32'h44e36498} /* (24, 6, 31) {real, imag} */,
  {32'h44297ff7, 32'hc3d00429} /* (24, 6, 30) {real, imag} */,
  {32'hc1df437e, 32'hc1be778e} /* (24, 6, 29) {real, imag} */,
  {32'hc33e3cb6, 32'hc1774d84} /* (24, 6, 28) {real, imag} */,
  {32'h4353fbe0, 32'hc305979f} /* (24, 6, 27) {real, imag} */,
  {32'h3fcc3b30, 32'hc315ff8a} /* (24, 6, 26) {real, imag} */,
  {32'h41b7afa4, 32'hc2a095a8} /* (24, 6, 25) {real, imag} */,
  {32'h40d961c8, 32'hc0891d64} /* (24, 6, 24) {real, imag} */,
  {32'hc2108e16, 32'hc237cbd8} /* (24, 6, 23) {real, imag} */,
  {32'hc20604dc, 32'hc16bfcec} /* (24, 6, 22) {real, imag} */,
  {32'h41032135, 32'h41f6fa0d} /* (24, 6, 21) {real, imag} */,
  {32'hc21de002, 32'h420bfa8a} /* (24, 6, 20) {real, imag} */,
  {32'h420b5fc0, 32'hc10b0ad6} /* (24, 6, 19) {real, imag} */,
  {32'h42599a0b, 32'hc252eac3} /* (24, 6, 18) {real, imag} */,
  {32'hc1bf6214, 32'h40ca4ef8} /* (24, 6, 17) {real, imag} */,
  {32'hbf9f3380, 32'h00000000} /* (24, 6, 16) {real, imag} */,
  {32'hc1bf6214, 32'hc0ca4ef8} /* (24, 6, 15) {real, imag} */,
  {32'h42599a0b, 32'h4252eac3} /* (24, 6, 14) {real, imag} */,
  {32'h420b5fc0, 32'h410b0ad6} /* (24, 6, 13) {real, imag} */,
  {32'hc21de002, 32'hc20bfa8a} /* (24, 6, 12) {real, imag} */,
  {32'h41032135, 32'hc1f6fa0d} /* (24, 6, 11) {real, imag} */,
  {32'hc20604dc, 32'h416bfcec} /* (24, 6, 10) {real, imag} */,
  {32'hc2108e16, 32'h4237cbd8} /* (24, 6, 9) {real, imag} */,
  {32'h40d961c8, 32'h40891d64} /* (24, 6, 8) {real, imag} */,
  {32'h41b7afa4, 32'h42a095a8} /* (24, 6, 7) {real, imag} */,
  {32'h3fcc3b30, 32'h4315ff8a} /* (24, 6, 6) {real, imag} */,
  {32'h4353fbe0, 32'h4305979f} /* (24, 6, 5) {real, imag} */,
  {32'hc33e3cb6, 32'h41774d84} /* (24, 6, 4) {real, imag} */,
  {32'hc1df437e, 32'h41be778e} /* (24, 6, 3) {real, imag} */,
  {32'h44297ff7, 32'h43d00429} /* (24, 6, 2) {real, imag} */,
  {32'hc52d7c4b, 32'hc4e36498} /* (24, 6, 1) {real, imag} */,
  {32'hc568ad58, 32'h00000000} /* (24, 6, 0) {real, imag} */,
  {32'hc529762e, 32'h4518d1a0} /* (24, 5, 31) {real, imag} */,
  {32'h4344db00, 32'hc40e0164} /* (24, 5, 30) {real, imag} */,
  {32'h4283a1b9, 32'h42ddfcda} /* (24, 5, 29) {real, imag} */,
  {32'h42482ec3, 32'hc2e16640} /* (24, 5, 28) {real, imag} */,
  {32'h42c92f2f, 32'h420600aa} /* (24, 5, 27) {real, imag} */,
  {32'h422cdf03, 32'hc2ab1632} /* (24, 5, 26) {real, imag} */,
  {32'h41e08bed, 32'h42c41014} /* (24, 5, 25) {real, imag} */,
  {32'hc1cc6c56, 32'hc2cf58b9} /* (24, 5, 24) {real, imag} */,
  {32'hc2a57ef7, 32'h424cb4b9} /* (24, 5, 23) {real, imag} */,
  {32'h404efe90, 32'hc12c5682} /* (24, 5, 22) {real, imag} */,
  {32'hc2906629, 32'h40d06462} /* (24, 5, 21) {real, imag} */,
  {32'hc13fc0f6, 32'hc236d0b0} /* (24, 5, 20) {real, imag} */,
  {32'h41d56f9a, 32'hc180284e} /* (24, 5, 19) {real, imag} */,
  {32'hc25eda3c, 32'hc24df555} /* (24, 5, 18) {real, imag} */,
  {32'h4165a7e9, 32'h41369d0e} /* (24, 5, 17) {real, imag} */,
  {32'h42c549e4, 32'h00000000} /* (24, 5, 16) {real, imag} */,
  {32'h4165a7e9, 32'hc1369d0e} /* (24, 5, 15) {real, imag} */,
  {32'hc25eda3c, 32'h424df555} /* (24, 5, 14) {real, imag} */,
  {32'h41d56f9a, 32'h4180284e} /* (24, 5, 13) {real, imag} */,
  {32'hc13fc0f6, 32'h4236d0b0} /* (24, 5, 12) {real, imag} */,
  {32'hc2906629, 32'hc0d06462} /* (24, 5, 11) {real, imag} */,
  {32'h404efe90, 32'h412c5682} /* (24, 5, 10) {real, imag} */,
  {32'hc2a57ef7, 32'hc24cb4b9} /* (24, 5, 9) {real, imag} */,
  {32'hc1cc6c56, 32'h42cf58b9} /* (24, 5, 8) {real, imag} */,
  {32'h41e08bed, 32'hc2c41014} /* (24, 5, 7) {real, imag} */,
  {32'h422cdf03, 32'h42ab1632} /* (24, 5, 6) {real, imag} */,
  {32'h42c92f2f, 32'hc20600aa} /* (24, 5, 5) {real, imag} */,
  {32'h42482ec3, 32'h42e16640} /* (24, 5, 4) {real, imag} */,
  {32'h4283a1b9, 32'hc2ddfcda} /* (24, 5, 3) {real, imag} */,
  {32'h4344db00, 32'h440e0164} /* (24, 5, 2) {real, imag} */,
  {32'hc529762e, 32'hc518d1a0} /* (24, 5, 1) {real, imag} */,
  {32'hc574b4a2, 32'h00000000} /* (24, 5, 0) {real, imag} */,
  {32'hc51be12b, 32'h45365fc3} /* (24, 4, 31) {real, imag} */,
  {32'hc33e7ff2, 32'hc42f99b4} /* (24, 4, 30) {real, imag} */,
  {32'h42438419, 32'h418f85d0} /* (24, 4, 29) {real, imag} */,
  {32'h431a6a40, 32'hc34a9325} /* (24, 4, 28) {real, imag} */,
  {32'h42d5d8d2, 32'h42f5190e} /* (24, 4, 27) {real, imag} */,
  {32'h419b5f3c, 32'hc2078d0a} /* (24, 4, 26) {real, imag} */,
  {32'h428b0a4c, 32'h429e76fd} /* (24, 4, 25) {real, imag} */,
  {32'hc0a9b418, 32'hc2aed402} /* (24, 4, 24) {real, imag} */,
  {32'h41821958, 32'h41c284d5} /* (24, 4, 23) {real, imag} */,
  {32'h41ee1007, 32'hc29e6c92} /* (24, 4, 22) {real, imag} */,
  {32'h425bac2f, 32'h42240a6f} /* (24, 4, 21) {real, imag} */,
  {32'hc25f6f48, 32'hc127c0d8} /* (24, 4, 20) {real, imag} */,
  {32'h4269104d, 32'hc20fac2a} /* (24, 4, 19) {real, imag} */,
  {32'hc1a6d41b, 32'hc190e688} /* (24, 4, 18) {real, imag} */,
  {32'h417fa104, 32'hc28946ec} /* (24, 4, 17) {real, imag} */,
  {32'hc1463f2e, 32'h00000000} /* (24, 4, 16) {real, imag} */,
  {32'h417fa104, 32'h428946ec} /* (24, 4, 15) {real, imag} */,
  {32'hc1a6d41b, 32'h4190e688} /* (24, 4, 14) {real, imag} */,
  {32'h4269104d, 32'h420fac2a} /* (24, 4, 13) {real, imag} */,
  {32'hc25f6f48, 32'h4127c0d8} /* (24, 4, 12) {real, imag} */,
  {32'h425bac2f, 32'hc2240a6f} /* (24, 4, 11) {real, imag} */,
  {32'h41ee1007, 32'h429e6c92} /* (24, 4, 10) {real, imag} */,
  {32'h41821958, 32'hc1c284d5} /* (24, 4, 9) {real, imag} */,
  {32'hc0a9b418, 32'h42aed402} /* (24, 4, 8) {real, imag} */,
  {32'h428b0a4c, 32'hc29e76fd} /* (24, 4, 7) {real, imag} */,
  {32'h419b5f3c, 32'h42078d0a} /* (24, 4, 6) {real, imag} */,
  {32'h42d5d8d2, 32'hc2f5190e} /* (24, 4, 5) {real, imag} */,
  {32'h431a6a40, 32'h434a9325} /* (24, 4, 4) {real, imag} */,
  {32'h42438419, 32'hc18f85d0} /* (24, 4, 3) {real, imag} */,
  {32'hc33e7ff2, 32'h442f99b4} /* (24, 4, 2) {real, imag} */,
  {32'hc51be12b, 32'hc5365fc3} /* (24, 4, 1) {real, imag} */,
  {32'hc5833a5b, 32'h00000000} /* (24, 4, 0) {real, imag} */,
  {32'hc5238008, 32'h453edb8f} /* (24, 3, 31) {real, imag} */,
  {32'hc35f5336, 32'hc4387f7e} /* (24, 3, 30) {real, imag} */,
  {32'h43281676, 32'h427b49ba} /* (24, 3, 29) {real, imag} */,
  {32'h430217c1, 32'hc36c8b05} /* (24, 3, 28) {real, imag} */,
  {32'h438b292f, 32'h42346cca} /* (24, 3, 27) {real, imag} */,
  {32'hc3094730, 32'hc219d18f} /* (24, 3, 26) {real, imag} */,
  {32'hc18b7cbe, 32'hc2a15589} /* (24, 3, 25) {real, imag} */,
  {32'hc2a67fa5, 32'hc17ddcf8} /* (24, 3, 24) {real, imag} */,
  {32'hc24e08a7, 32'hc19d3b29} /* (24, 3, 23) {real, imag} */,
  {32'h42bc324c, 32'hc27a29f0} /* (24, 3, 22) {real, imag} */,
  {32'h42a5192e, 32'h4193b07e} /* (24, 3, 21) {real, imag} */,
  {32'hbf40d380, 32'hc1c8cecb} /* (24, 3, 20) {real, imag} */,
  {32'h42418abf, 32'h42ab122c} /* (24, 3, 19) {real, imag} */,
  {32'h4114f4f8, 32'h41efb27a} /* (24, 3, 18) {real, imag} */,
  {32'h41200f5e, 32'hc206d758} /* (24, 3, 17) {real, imag} */,
  {32'hc22a9c5a, 32'h00000000} /* (24, 3, 16) {real, imag} */,
  {32'h41200f5e, 32'h4206d758} /* (24, 3, 15) {real, imag} */,
  {32'h4114f4f8, 32'hc1efb27a} /* (24, 3, 14) {real, imag} */,
  {32'h42418abf, 32'hc2ab122c} /* (24, 3, 13) {real, imag} */,
  {32'hbf40d380, 32'h41c8cecb} /* (24, 3, 12) {real, imag} */,
  {32'h42a5192e, 32'hc193b07e} /* (24, 3, 11) {real, imag} */,
  {32'h42bc324c, 32'h427a29f0} /* (24, 3, 10) {real, imag} */,
  {32'hc24e08a7, 32'h419d3b29} /* (24, 3, 9) {real, imag} */,
  {32'hc2a67fa5, 32'h417ddcf8} /* (24, 3, 8) {real, imag} */,
  {32'hc18b7cbe, 32'h42a15589} /* (24, 3, 7) {real, imag} */,
  {32'hc3094730, 32'h4219d18f} /* (24, 3, 6) {real, imag} */,
  {32'h438b292f, 32'hc2346cca} /* (24, 3, 5) {real, imag} */,
  {32'h430217c1, 32'h436c8b05} /* (24, 3, 4) {real, imag} */,
  {32'h43281676, 32'hc27b49ba} /* (24, 3, 3) {real, imag} */,
  {32'hc35f5336, 32'h44387f7e} /* (24, 3, 2) {real, imag} */,
  {32'hc5238008, 32'hc53edb8f} /* (24, 3, 1) {real, imag} */,
  {32'hc582a3e5, 32'h00000000} /* (24, 3, 0) {real, imag} */,
  {32'hc51b7da7, 32'h4540b43a} /* (24, 2, 31) {real, imag} */,
  {32'hc3aad732, 32'hc43c44ed} /* (24, 2, 30) {real, imag} */,
  {32'h437366df, 32'h424b66f0} /* (24, 2, 29) {real, imag} */,
  {32'h42d67e20, 32'hc3987288} /* (24, 2, 28) {real, imag} */,
  {32'h43062c0e, 32'hbec24480} /* (24, 2, 27) {real, imag} */,
  {32'h42621a5d, 32'h426a50ec} /* (24, 2, 26) {real, imag} */,
  {32'hc13ed094, 32'h422de2ba} /* (24, 2, 25) {real, imag} */,
  {32'h41b19444, 32'h423a73e2} /* (24, 2, 24) {real, imag} */,
  {32'hc20e006a, 32'hc1f3e03a} /* (24, 2, 23) {real, imag} */,
  {32'h42823ff8, 32'hc2a2f2bc} /* (24, 2, 22) {real, imag} */,
  {32'h4240bbd9, 32'h3f384200} /* (24, 2, 21) {real, imag} */,
  {32'hc28c6d56, 32'hc2aa61ed} /* (24, 2, 20) {real, imag} */,
  {32'h428c5d05, 32'h41299172} /* (24, 2, 19) {real, imag} */,
  {32'hc1f5eebe, 32'h41d49d58} /* (24, 2, 18) {real, imag} */,
  {32'hc21e84d6, 32'h41b4dd0c} /* (24, 2, 17) {real, imag} */,
  {32'h41a0a15c, 32'h00000000} /* (24, 2, 16) {real, imag} */,
  {32'hc21e84d6, 32'hc1b4dd0c} /* (24, 2, 15) {real, imag} */,
  {32'hc1f5eebe, 32'hc1d49d58} /* (24, 2, 14) {real, imag} */,
  {32'h428c5d05, 32'hc1299172} /* (24, 2, 13) {real, imag} */,
  {32'hc28c6d56, 32'h42aa61ed} /* (24, 2, 12) {real, imag} */,
  {32'h4240bbd9, 32'hbf384200} /* (24, 2, 11) {real, imag} */,
  {32'h42823ff8, 32'h42a2f2bc} /* (24, 2, 10) {real, imag} */,
  {32'hc20e006a, 32'h41f3e03a} /* (24, 2, 9) {real, imag} */,
  {32'h41b19444, 32'hc23a73e2} /* (24, 2, 8) {real, imag} */,
  {32'hc13ed094, 32'hc22de2ba} /* (24, 2, 7) {real, imag} */,
  {32'h42621a5d, 32'hc26a50ec} /* (24, 2, 6) {real, imag} */,
  {32'h43062c0e, 32'h3ec24480} /* (24, 2, 5) {real, imag} */,
  {32'h42d67e20, 32'h43987288} /* (24, 2, 4) {real, imag} */,
  {32'h437366df, 32'hc24b66f0} /* (24, 2, 3) {real, imag} */,
  {32'hc3aad732, 32'h443c44ed} /* (24, 2, 2) {real, imag} */,
  {32'hc51b7da7, 32'hc540b43a} /* (24, 2, 1) {real, imag} */,
  {32'hc5822409, 32'h00000000} /* (24, 2, 0) {real, imag} */,
  {32'hc5226249, 32'h45307d30} /* (24, 1, 31) {real, imag} */,
  {32'hc31e8a3a, 32'hc421ecfd} /* (24, 1, 30) {real, imag} */,
  {32'h4386286e, 32'hbd3cb500} /* (24, 1, 29) {real, imag} */,
  {32'h432f59be, 32'hc38a8ae6} /* (24, 1, 28) {real, imag} */,
  {32'h42ab3f0f, 32'h4128539e} /* (24, 1, 27) {real, imag} */,
  {32'h41dcb41e, 32'hc25cffea} /* (24, 1, 26) {real, imag} */,
  {32'hc28cf9e0, 32'h42a427ca} /* (24, 1, 25) {real, imag} */,
  {32'h421cd6d2, 32'hc284e8a2} /* (24, 1, 24) {real, imag} */,
  {32'h4216ece6, 32'hc1c7340f} /* (24, 1, 23) {real, imag} */,
  {32'hc184cd0a, 32'h4201762e} /* (24, 1, 22) {real, imag} */,
  {32'h40f04446, 32'hc2017486} /* (24, 1, 21) {real, imag} */,
  {32'hc221dec0, 32'h41e3c560} /* (24, 1, 20) {real, imag} */,
  {32'hc10541b0, 32'h4224ac5f} /* (24, 1, 19) {real, imag} */,
  {32'h418700c8, 32'hc2aba606} /* (24, 1, 18) {real, imag} */,
  {32'h41a79a98, 32'h42ba9d8f} /* (24, 1, 17) {real, imag} */,
  {32'h4214b840, 32'h00000000} /* (24, 1, 16) {real, imag} */,
  {32'h41a79a98, 32'hc2ba9d8f} /* (24, 1, 15) {real, imag} */,
  {32'h418700c8, 32'h42aba606} /* (24, 1, 14) {real, imag} */,
  {32'hc10541b0, 32'hc224ac5f} /* (24, 1, 13) {real, imag} */,
  {32'hc221dec0, 32'hc1e3c560} /* (24, 1, 12) {real, imag} */,
  {32'h40f04446, 32'h42017486} /* (24, 1, 11) {real, imag} */,
  {32'hc184cd0a, 32'hc201762e} /* (24, 1, 10) {real, imag} */,
  {32'h4216ece6, 32'h41c7340f} /* (24, 1, 9) {real, imag} */,
  {32'h421cd6d2, 32'h4284e8a2} /* (24, 1, 8) {real, imag} */,
  {32'hc28cf9e0, 32'hc2a427ca} /* (24, 1, 7) {real, imag} */,
  {32'h41dcb41e, 32'h425cffea} /* (24, 1, 6) {real, imag} */,
  {32'h42ab3f0f, 32'hc128539e} /* (24, 1, 5) {real, imag} */,
  {32'h432f59be, 32'h438a8ae6} /* (24, 1, 4) {real, imag} */,
  {32'h4386286e, 32'h3d3cb500} /* (24, 1, 3) {real, imag} */,
  {32'hc31e8a3a, 32'h4421ecfd} /* (24, 1, 2) {real, imag} */,
  {32'hc5226249, 32'hc5307d30} /* (24, 1, 1) {real, imag} */,
  {32'hc582bb5c, 32'h00000000} /* (24, 1, 0) {real, imag} */,
  {32'hc52de981, 32'h450b29c4} /* (24, 0, 31) {real, imag} */,
  {32'h42e7727c, 32'hc39a0146} /* (24, 0, 30) {real, imag} */,
  {32'h432e5ae1, 32'hc16b19f6} /* (24, 0, 29) {real, imag} */,
  {32'h42dfdf48, 32'hc318cb4e} /* (24, 0, 28) {real, imag} */,
  {32'h42bb7a74, 32'h41b839ad} /* (24, 0, 27) {real, imag} */,
  {32'hc20d0566, 32'hc1300c6e} /* (24, 0, 26) {real, imag} */,
  {32'hc1835108, 32'hc1149e6e} /* (24, 0, 25) {real, imag} */,
  {32'h419f58a8, 32'h410c63c8} /* (24, 0, 24) {real, imag} */,
  {32'h42824eb6, 32'hc1ea97bc} /* (24, 0, 23) {real, imag} */,
  {32'hc2c26272, 32'hc10f9be4} /* (24, 0, 22) {real, imag} */,
  {32'h40c65739, 32'hc1ded516} /* (24, 0, 21) {real, imag} */,
  {32'h405bcb92, 32'h41d630cd} /* (24, 0, 20) {real, imag} */,
  {32'h40d7a88e, 32'h420a2924} /* (24, 0, 19) {real, imag} */,
  {32'hc14b34b7, 32'hc0c04b2a} /* (24, 0, 18) {real, imag} */,
  {32'hc21c984d, 32'hc0ed79ec} /* (24, 0, 17) {real, imag} */,
  {32'h422190b2, 32'h00000000} /* (24, 0, 16) {real, imag} */,
  {32'hc21c984d, 32'h40ed79ec} /* (24, 0, 15) {real, imag} */,
  {32'hc14b34b7, 32'h40c04b2a} /* (24, 0, 14) {real, imag} */,
  {32'h40d7a88e, 32'hc20a2924} /* (24, 0, 13) {real, imag} */,
  {32'h405bcb92, 32'hc1d630cd} /* (24, 0, 12) {real, imag} */,
  {32'h40c65739, 32'h41ded516} /* (24, 0, 11) {real, imag} */,
  {32'hc2c26272, 32'h410f9be4} /* (24, 0, 10) {real, imag} */,
  {32'h42824eb6, 32'h41ea97bc} /* (24, 0, 9) {real, imag} */,
  {32'h419f58a8, 32'hc10c63c8} /* (24, 0, 8) {real, imag} */,
  {32'hc1835108, 32'h41149e6e} /* (24, 0, 7) {real, imag} */,
  {32'hc20d0566, 32'h41300c6e} /* (24, 0, 6) {real, imag} */,
  {32'h42bb7a74, 32'hc1b839ad} /* (24, 0, 5) {real, imag} */,
  {32'h42dfdf48, 32'h4318cb4e} /* (24, 0, 4) {real, imag} */,
  {32'h432e5ae1, 32'h416b19f6} /* (24, 0, 3) {real, imag} */,
  {32'h42e7727c, 32'h439a0146} /* (24, 0, 2) {real, imag} */,
  {32'hc52de981, 32'hc50b29c4} /* (24, 0, 1) {real, imag} */,
  {32'hc580ece3, 32'h00000000} /* (24, 0, 0) {real, imag} */,
  {32'hc567ece0, 32'h45048bc6} /* (23, 31, 31) {real, imag} */,
  {32'h4434a48c, 32'hc3a15588} /* (23, 31, 30) {real, imag} */,
  {32'h4285f1cd, 32'h412b7f4a} /* (23, 31, 29) {real, imag} */,
  {32'hc2de2430, 32'hc18e2e40} /* (23, 31, 28) {real, imag} */,
  {32'h42fb60a4, 32'h410f0c06} /* (23, 31, 27) {real, imag} */,
  {32'h404cc460, 32'h42251112} /* (23, 31, 26) {real, imag} */,
  {32'hc2220f2c, 32'h428f8000} /* (23, 31, 25) {real, imag} */,
  {32'h42befa4f, 32'hc236c5ca} /* (23, 31, 24) {real, imag} */,
  {32'hc01e2440, 32'hc2f13846} /* (23, 31, 23) {real, imag} */,
  {32'hc234127e, 32'h42896780} /* (23, 31, 22) {real, imag} */,
  {32'h42393498, 32'h40fde72c} /* (23, 31, 21) {real, imag} */,
  {32'hc25ffae4, 32'hc1da5f19} /* (23, 31, 20) {real, imag} */,
  {32'h42192f2e, 32'hc1597fb1} /* (23, 31, 19) {real, imag} */,
  {32'h421d7fb8, 32'hc261bdc7} /* (23, 31, 18) {real, imag} */,
  {32'hc12a9538, 32'h40b7dd0c} /* (23, 31, 17) {real, imag} */,
  {32'hc28bf111, 32'h00000000} /* (23, 31, 16) {real, imag} */,
  {32'hc12a9538, 32'hc0b7dd0c} /* (23, 31, 15) {real, imag} */,
  {32'h421d7fb8, 32'h4261bdc7} /* (23, 31, 14) {real, imag} */,
  {32'h42192f2e, 32'h41597fb1} /* (23, 31, 13) {real, imag} */,
  {32'hc25ffae4, 32'h41da5f19} /* (23, 31, 12) {real, imag} */,
  {32'h42393498, 32'hc0fde72c} /* (23, 31, 11) {real, imag} */,
  {32'hc234127e, 32'hc2896780} /* (23, 31, 10) {real, imag} */,
  {32'hc01e2440, 32'h42f13846} /* (23, 31, 9) {real, imag} */,
  {32'h42befa4f, 32'h4236c5ca} /* (23, 31, 8) {real, imag} */,
  {32'hc2220f2c, 32'hc28f8000} /* (23, 31, 7) {real, imag} */,
  {32'h404cc460, 32'hc2251112} /* (23, 31, 6) {real, imag} */,
  {32'h42fb60a4, 32'hc10f0c06} /* (23, 31, 5) {real, imag} */,
  {32'hc2de2430, 32'h418e2e40} /* (23, 31, 4) {real, imag} */,
  {32'h4285f1cd, 32'hc12b7f4a} /* (23, 31, 3) {real, imag} */,
  {32'h4434a48c, 32'h43a15588} /* (23, 31, 2) {real, imag} */,
  {32'hc567ece0, 32'hc5048bc6} /* (23, 31, 1) {real, imag} */,
  {32'hc597c953, 32'h00000000} /* (23, 31, 0) {real, imag} */,
  {32'hc582658f, 32'h44e7d93c} /* (23, 30, 31) {real, imag} */,
  {32'h448ed35d, 32'hc399c8b5} /* (23, 30, 30) {real, imag} */,
  {32'h42402462, 32'hc2427d0c} /* (23, 30, 29) {real, imag} */,
  {32'hc339d63e, 32'h42a0cae8} /* (23, 30, 28) {real, imag} */,
  {32'h4353f456, 32'hc2b50f5f} /* (23, 30, 27) {real, imag} */,
  {32'h43227f6b, 32'h42b35a1e} /* (23, 30, 26) {real, imag} */,
  {32'hc31749aa, 32'h4279d960} /* (23, 30, 25) {real, imag} */,
  {32'h42633ca5, 32'hc2d52212} /* (23, 30, 24) {real, imag} */,
  {32'h420738fe, 32'h4127d9cc} /* (23, 30, 23) {real, imag} */,
  {32'hc142185e, 32'h423af091} /* (23, 30, 22) {real, imag} */,
  {32'hc28b33f3, 32'hc305b733} /* (23, 30, 21) {real, imag} */,
  {32'hc2a32415, 32'hc0dd2c70} /* (23, 30, 20) {real, imag} */,
  {32'hc1dfc1f9, 32'h421f08d4} /* (23, 30, 19) {real, imag} */,
  {32'h42a827fc, 32'hc2908115} /* (23, 30, 18) {real, imag} */,
  {32'hc25f0f05, 32'h4260ed0c} /* (23, 30, 17) {real, imag} */,
  {32'h41e3418f, 32'h00000000} /* (23, 30, 16) {real, imag} */,
  {32'hc25f0f05, 32'hc260ed0c} /* (23, 30, 15) {real, imag} */,
  {32'h42a827fc, 32'h42908115} /* (23, 30, 14) {real, imag} */,
  {32'hc1dfc1f9, 32'hc21f08d4} /* (23, 30, 13) {real, imag} */,
  {32'hc2a32415, 32'h40dd2c70} /* (23, 30, 12) {real, imag} */,
  {32'hc28b33f3, 32'h4305b733} /* (23, 30, 11) {real, imag} */,
  {32'hc142185e, 32'hc23af091} /* (23, 30, 10) {real, imag} */,
  {32'h420738fe, 32'hc127d9cc} /* (23, 30, 9) {real, imag} */,
  {32'h42633ca5, 32'h42d52212} /* (23, 30, 8) {real, imag} */,
  {32'hc31749aa, 32'hc279d960} /* (23, 30, 7) {real, imag} */,
  {32'h43227f6b, 32'hc2b35a1e} /* (23, 30, 6) {real, imag} */,
  {32'h4353f456, 32'h42b50f5f} /* (23, 30, 5) {real, imag} */,
  {32'hc339d63e, 32'hc2a0cae8} /* (23, 30, 4) {real, imag} */,
  {32'h42402462, 32'h42427d0c} /* (23, 30, 3) {real, imag} */,
  {32'h448ed35d, 32'h4399c8b5} /* (23, 30, 2) {real, imag} */,
  {32'hc582658f, 32'hc4e7d93c} /* (23, 30, 1) {real, imag} */,
  {32'hc59d1de8, 32'h00000000} /* (23, 30, 0) {real, imag} */,
  {32'hc58b4758, 32'h44c3c435} /* (23, 29, 31) {real, imag} */,
  {32'h44ae2864, 32'hc36bcb24} /* (23, 29, 30) {real, imag} */,
  {32'hc15ceb8c, 32'hc2c48813} /* (23, 29, 29) {real, imag} */,
  {32'hc370269a, 32'h43020bc6} /* (23, 29, 28) {real, imag} */,
  {32'h42077f44, 32'hc34601d3} /* (23, 29, 27) {real, imag} */,
  {32'h42a90076, 32'h423cf0d5} /* (23, 29, 26) {real, imag} */,
  {32'h420ed871, 32'hc19828d0} /* (23, 29, 25) {real, imag} */,
  {32'hc2073735, 32'hc2c66296} /* (23, 29, 24) {real, imag} */,
  {32'h41e0c00c, 32'h3ed5e4c0} /* (23, 29, 23) {real, imag} */,
  {32'h4285f6e2, 32'h3f72c780} /* (23, 29, 22) {real, imag} */,
  {32'h425cbec2, 32'hc0945920} /* (23, 29, 21) {real, imag} */,
  {32'h42541214, 32'hc15a93ed} /* (23, 29, 20) {real, imag} */,
  {32'h41b4c05c, 32'hc1793432} /* (23, 29, 19) {real, imag} */,
  {32'hc28d70b6, 32'h41118948} /* (23, 29, 18) {real, imag} */,
  {32'hc1acc649, 32'h408e2e8c} /* (23, 29, 17) {real, imag} */,
  {32'h41cfb844, 32'h00000000} /* (23, 29, 16) {real, imag} */,
  {32'hc1acc649, 32'hc08e2e8c} /* (23, 29, 15) {real, imag} */,
  {32'hc28d70b6, 32'hc1118948} /* (23, 29, 14) {real, imag} */,
  {32'h41b4c05c, 32'h41793432} /* (23, 29, 13) {real, imag} */,
  {32'h42541214, 32'h415a93ed} /* (23, 29, 12) {real, imag} */,
  {32'h425cbec2, 32'h40945920} /* (23, 29, 11) {real, imag} */,
  {32'h4285f6e2, 32'hbf72c780} /* (23, 29, 10) {real, imag} */,
  {32'h41e0c00c, 32'hbed5e4c0} /* (23, 29, 9) {real, imag} */,
  {32'hc2073735, 32'h42c66296} /* (23, 29, 8) {real, imag} */,
  {32'h420ed871, 32'h419828d0} /* (23, 29, 7) {real, imag} */,
  {32'h42a90076, 32'hc23cf0d5} /* (23, 29, 6) {real, imag} */,
  {32'h42077f44, 32'h434601d3} /* (23, 29, 5) {real, imag} */,
  {32'hc370269a, 32'hc3020bc6} /* (23, 29, 4) {real, imag} */,
  {32'hc15ceb8c, 32'h42c48813} /* (23, 29, 3) {real, imag} */,
  {32'h44ae2864, 32'h436bcb24} /* (23, 29, 2) {real, imag} */,
  {32'hc58b4758, 32'hc4c3c435} /* (23, 29, 1) {real, imag} */,
  {32'hc5a06884, 32'h00000000} /* (23, 29, 0) {real, imag} */,
  {32'hc593ead0, 32'h4498881e} /* (23, 28, 31) {real, imag} */,
  {32'h44c15bd9, 32'hc39826e8} /* (23, 28, 30) {real, imag} */,
  {32'hc244152e, 32'hc1f9c5b8} /* (23, 28, 29) {real, imag} */,
  {32'hc379b573, 32'h429ac417} /* (23, 28, 28) {real, imag} */,
  {32'h42bb3438, 32'hc2dc065b} /* (23, 28, 27) {real, imag} */,
  {32'h430e3a69, 32'hc0906d18} /* (23, 28, 26) {real, imag} */,
  {32'h42a80e50, 32'h42beb484} /* (23, 28, 25) {real, imag} */,
  {32'h4254379a, 32'hc27a47aa} /* (23, 28, 24) {real, imag} */,
  {32'hc0b037f8, 32'h429ad6ee} /* (23, 28, 23) {real, imag} */,
  {32'h429a02c5, 32'h42467cf0} /* (23, 28, 22) {real, imag} */,
  {32'h42b84883, 32'h42030d86} /* (23, 28, 21) {real, imag} */,
  {32'hc1cf41de, 32'h41bf1776} /* (23, 28, 20) {real, imag} */,
  {32'h41319dff, 32'hc20306a8} /* (23, 28, 19) {real, imag} */,
  {32'h423d9de1, 32'h41c9b820} /* (23, 28, 18) {real, imag} */,
  {32'h4230faa5, 32'h42361330} /* (23, 28, 17) {real, imag} */,
  {32'h4263a37a, 32'h00000000} /* (23, 28, 16) {real, imag} */,
  {32'h4230faa5, 32'hc2361330} /* (23, 28, 15) {real, imag} */,
  {32'h423d9de1, 32'hc1c9b820} /* (23, 28, 14) {real, imag} */,
  {32'h41319dff, 32'h420306a8} /* (23, 28, 13) {real, imag} */,
  {32'hc1cf41de, 32'hc1bf1776} /* (23, 28, 12) {real, imag} */,
  {32'h42b84883, 32'hc2030d86} /* (23, 28, 11) {real, imag} */,
  {32'h429a02c5, 32'hc2467cf0} /* (23, 28, 10) {real, imag} */,
  {32'hc0b037f8, 32'hc29ad6ee} /* (23, 28, 9) {real, imag} */,
  {32'h4254379a, 32'h427a47aa} /* (23, 28, 8) {real, imag} */,
  {32'h42a80e50, 32'hc2beb484} /* (23, 28, 7) {real, imag} */,
  {32'h430e3a69, 32'h40906d18} /* (23, 28, 6) {real, imag} */,
  {32'h42bb3438, 32'h42dc065b} /* (23, 28, 5) {real, imag} */,
  {32'hc379b573, 32'hc29ac417} /* (23, 28, 4) {real, imag} */,
  {32'hc244152e, 32'h41f9c5b8} /* (23, 28, 3) {real, imag} */,
  {32'h44c15bd9, 32'h439826e8} /* (23, 28, 2) {real, imag} */,
  {32'hc593ead0, 32'hc498881e} /* (23, 28, 1) {real, imag} */,
  {32'hc5a223d2, 32'h00000000} /* (23, 28, 0) {real, imag} */,
  {32'hc593c2ba, 32'h44801ee0} /* (23, 27, 31) {real, imag} */,
  {32'h44c514ae, 32'hc37ffa10} /* (23, 27, 30) {real, imag} */,
  {32'h42e5aeb6, 32'hc264a0ac} /* (23, 27, 29) {real, imag} */,
  {32'hc29290e6, 32'h41d47ace} /* (23, 27, 28) {real, imag} */,
  {32'h43674efc, 32'hc330a882} /* (23, 27, 27) {real, imag} */,
  {32'h4280a7b7, 32'h43152c42} /* (23, 27, 26) {real, imag} */,
  {32'h424591ec, 32'h42851dc6} /* (23, 27, 25) {real, imag} */,
  {32'h428337e6, 32'h4118944d} /* (23, 27, 24) {real, imag} */,
  {32'h429a67cc, 32'h42afe520} /* (23, 27, 23) {real, imag} */,
  {32'h411820c4, 32'h40761420} /* (23, 27, 22) {real, imag} */,
  {32'hc2383d02, 32'hc28f7858} /* (23, 27, 21) {real, imag} */,
  {32'hc1241407, 32'hc22c238b} /* (23, 27, 20) {real, imag} */,
  {32'hc2f11411, 32'h41af8864} /* (23, 27, 19) {real, imag} */,
  {32'hc23557c8, 32'hc25a7a38} /* (23, 27, 18) {real, imag} */,
  {32'hc204e68e, 32'hc08fc420} /* (23, 27, 17) {real, imag} */,
  {32'hc1549e34, 32'h00000000} /* (23, 27, 16) {real, imag} */,
  {32'hc204e68e, 32'h408fc420} /* (23, 27, 15) {real, imag} */,
  {32'hc23557c8, 32'h425a7a38} /* (23, 27, 14) {real, imag} */,
  {32'hc2f11411, 32'hc1af8864} /* (23, 27, 13) {real, imag} */,
  {32'hc1241407, 32'h422c238b} /* (23, 27, 12) {real, imag} */,
  {32'hc2383d02, 32'h428f7858} /* (23, 27, 11) {real, imag} */,
  {32'h411820c4, 32'hc0761420} /* (23, 27, 10) {real, imag} */,
  {32'h429a67cc, 32'hc2afe520} /* (23, 27, 9) {real, imag} */,
  {32'h428337e6, 32'hc118944d} /* (23, 27, 8) {real, imag} */,
  {32'h424591ec, 32'hc2851dc6} /* (23, 27, 7) {real, imag} */,
  {32'h4280a7b7, 32'hc3152c42} /* (23, 27, 6) {real, imag} */,
  {32'h43674efc, 32'h4330a882} /* (23, 27, 5) {real, imag} */,
  {32'hc29290e6, 32'hc1d47ace} /* (23, 27, 4) {real, imag} */,
  {32'h42e5aeb6, 32'h4264a0ac} /* (23, 27, 3) {real, imag} */,
  {32'h44c514ae, 32'h437ffa10} /* (23, 27, 2) {real, imag} */,
  {32'hc593c2ba, 32'hc4801ee0} /* (23, 27, 1) {real, imag} */,
  {32'hc5a3565d, 32'h00000000} /* (23, 27, 0) {real, imag} */,
  {32'hc58d02b3, 32'h447407d1} /* (23, 26, 31) {real, imag} */,
  {32'h44caa5ec, 32'hc299891c} /* (23, 26, 30) {real, imag} */,
  {32'h428f5127, 32'hc2be0df0} /* (23, 26, 29) {real, imag} */,
  {32'hc2fbc75e, 32'hc06a5130} /* (23, 26, 28) {real, imag} */,
  {32'h431a5345, 32'hc33612aa} /* (23, 26, 27) {real, imag} */,
  {32'hc1919a36, 32'hc02015f8} /* (23, 26, 26) {real, imag} */,
  {32'hc1147398, 32'h4285d61f} /* (23, 26, 25) {real, imag} */,
  {32'h41d2995a, 32'h41d7d419} /* (23, 26, 24) {real, imag} */,
  {32'h42ba969c, 32'hc1c39fa1} /* (23, 26, 23) {real, imag} */,
  {32'hc30a5c64, 32'hc257c656} /* (23, 26, 22) {real, imag} */,
  {32'h41d549ae, 32'h41891b1e} /* (23, 26, 21) {real, imag} */,
  {32'h4143a2cc, 32'h41922d72} /* (23, 26, 20) {real, imag} */,
  {32'h4240a0a0, 32'h4209a8b0} /* (23, 26, 19) {real, imag} */,
  {32'hc206fb68, 32'h41d08419} /* (23, 26, 18) {real, imag} */,
  {32'h411f49e2, 32'hc187b1e4} /* (23, 26, 17) {real, imag} */,
  {32'hc2b57969, 32'h00000000} /* (23, 26, 16) {real, imag} */,
  {32'h411f49e2, 32'h4187b1e4} /* (23, 26, 15) {real, imag} */,
  {32'hc206fb68, 32'hc1d08419} /* (23, 26, 14) {real, imag} */,
  {32'h4240a0a0, 32'hc209a8b0} /* (23, 26, 13) {real, imag} */,
  {32'h4143a2cc, 32'hc1922d72} /* (23, 26, 12) {real, imag} */,
  {32'h41d549ae, 32'hc1891b1e} /* (23, 26, 11) {real, imag} */,
  {32'hc30a5c64, 32'h4257c656} /* (23, 26, 10) {real, imag} */,
  {32'h42ba969c, 32'h41c39fa1} /* (23, 26, 9) {real, imag} */,
  {32'h41d2995a, 32'hc1d7d419} /* (23, 26, 8) {real, imag} */,
  {32'hc1147398, 32'hc285d61f} /* (23, 26, 7) {real, imag} */,
  {32'hc1919a36, 32'h402015f8} /* (23, 26, 6) {real, imag} */,
  {32'h431a5345, 32'h433612aa} /* (23, 26, 5) {real, imag} */,
  {32'hc2fbc75e, 32'h406a5130} /* (23, 26, 4) {real, imag} */,
  {32'h428f5127, 32'h42be0df0} /* (23, 26, 3) {real, imag} */,
  {32'h44caa5ec, 32'h4299891c} /* (23, 26, 2) {real, imag} */,
  {32'hc58d02b3, 32'hc47407d1} /* (23, 26, 1) {real, imag} */,
  {32'hc59cf28f, 32'h00000000} /* (23, 26, 0) {real, imag} */,
  {32'hc586d72f, 32'h44338da9} /* (23, 25, 31) {real, imag} */,
  {32'h44cdbaf4, 32'hc30bafb0} /* (23, 25, 30) {real, imag} */,
  {32'hc227de3c, 32'h40649950} /* (23, 25, 29) {real, imag} */,
  {32'hc30fe36c, 32'hc1de198a} /* (23, 25, 28) {real, imag} */,
  {32'h43af554b, 32'h4070a6c0} /* (23, 25, 27) {real, imag} */,
  {32'h41da70c3, 32'h429bbeb6} /* (23, 25, 26) {real, imag} */,
  {32'h42cd90f2, 32'hc099606c} /* (23, 25, 25) {real, imag} */,
  {32'h430d2452, 32'hc1be49e8} /* (23, 25, 24) {real, imag} */,
  {32'h41758f0c, 32'h4297837a} /* (23, 25, 23) {real, imag} */,
  {32'hc0f0ce6a, 32'h4209d626} /* (23, 25, 22) {real, imag} */,
  {32'h421b6bdd, 32'hc28a201f} /* (23, 25, 21) {real, imag} */,
  {32'h4262def9, 32'h41e98330} /* (23, 25, 20) {real, imag} */,
  {32'hc11a8f74, 32'h408e0b38} /* (23, 25, 19) {real, imag} */,
  {32'hc101fbc0, 32'hc2258fa9} /* (23, 25, 18) {real, imag} */,
  {32'hc136457e, 32'h427fa26d} /* (23, 25, 17) {real, imag} */,
  {32'hc1f9214d, 32'h00000000} /* (23, 25, 16) {real, imag} */,
  {32'hc136457e, 32'hc27fa26d} /* (23, 25, 15) {real, imag} */,
  {32'hc101fbc0, 32'h42258fa9} /* (23, 25, 14) {real, imag} */,
  {32'hc11a8f74, 32'hc08e0b38} /* (23, 25, 13) {real, imag} */,
  {32'h4262def9, 32'hc1e98330} /* (23, 25, 12) {real, imag} */,
  {32'h421b6bdd, 32'h428a201f} /* (23, 25, 11) {real, imag} */,
  {32'hc0f0ce6a, 32'hc209d626} /* (23, 25, 10) {real, imag} */,
  {32'h41758f0c, 32'hc297837a} /* (23, 25, 9) {real, imag} */,
  {32'h430d2452, 32'h41be49e8} /* (23, 25, 8) {real, imag} */,
  {32'h42cd90f2, 32'h4099606c} /* (23, 25, 7) {real, imag} */,
  {32'h41da70c3, 32'hc29bbeb6} /* (23, 25, 6) {real, imag} */,
  {32'h43af554b, 32'hc070a6c0} /* (23, 25, 5) {real, imag} */,
  {32'hc30fe36c, 32'h41de198a} /* (23, 25, 4) {real, imag} */,
  {32'hc227de3c, 32'hc0649950} /* (23, 25, 3) {real, imag} */,
  {32'h44cdbaf4, 32'h430bafb0} /* (23, 25, 2) {real, imag} */,
  {32'hc586d72f, 32'hc4338da9} /* (23, 25, 1) {real, imag} */,
  {32'hc58faa32, 32'h00000000} /* (23, 25, 0) {real, imag} */,
  {32'hc57400dc, 32'h4402142f} /* (23, 24, 31) {real, imag} */,
  {32'h44c3bc78, 32'hc355a464} /* (23, 24, 30) {real, imag} */,
  {32'hc2b62828, 32'h42cbbfa6} /* (23, 24, 29) {real, imag} */,
  {32'hc1f6c75a, 32'h42054718} /* (23, 24, 28) {real, imag} */,
  {32'h43707912, 32'hc31c2b1a} /* (23, 24, 27) {real, imag} */,
  {32'h41041bc4, 32'hc2ad373c} /* (23, 24, 26) {real, imag} */,
  {32'h4241c535, 32'h41709520} /* (23, 24, 25) {real, imag} */,
  {32'h424e1bc0, 32'h42c99814} /* (23, 24, 24) {real, imag} */,
  {32'h41e2445a, 32'hc150d438} /* (23, 24, 23) {real, imag} */,
  {32'hc18f8319, 32'h42a44ce2} /* (23, 24, 22) {real, imag} */,
  {32'h42461941, 32'hc29aec9b} /* (23, 24, 21) {real, imag} */,
  {32'hc15b9a30, 32'h41b5308c} /* (23, 24, 20) {real, imag} */,
  {32'hc28b682c, 32'hc225e327} /* (23, 24, 19) {real, imag} */,
  {32'h41234bd4, 32'h422f62fb} /* (23, 24, 18) {real, imag} */,
  {32'hc1a3322a, 32'hc1b8abe4} /* (23, 24, 17) {real, imag} */,
  {32'h43037f4d, 32'h00000000} /* (23, 24, 16) {real, imag} */,
  {32'hc1a3322a, 32'h41b8abe4} /* (23, 24, 15) {real, imag} */,
  {32'h41234bd4, 32'hc22f62fb} /* (23, 24, 14) {real, imag} */,
  {32'hc28b682c, 32'h4225e327} /* (23, 24, 13) {real, imag} */,
  {32'hc15b9a30, 32'hc1b5308c} /* (23, 24, 12) {real, imag} */,
  {32'h42461941, 32'h429aec9b} /* (23, 24, 11) {real, imag} */,
  {32'hc18f8319, 32'hc2a44ce2} /* (23, 24, 10) {real, imag} */,
  {32'h41e2445a, 32'h4150d438} /* (23, 24, 9) {real, imag} */,
  {32'h424e1bc0, 32'hc2c99814} /* (23, 24, 8) {real, imag} */,
  {32'h4241c535, 32'hc1709520} /* (23, 24, 7) {real, imag} */,
  {32'h41041bc4, 32'h42ad373c} /* (23, 24, 6) {real, imag} */,
  {32'h43707912, 32'h431c2b1a} /* (23, 24, 5) {real, imag} */,
  {32'hc1f6c75a, 32'hc2054718} /* (23, 24, 4) {real, imag} */,
  {32'hc2b62828, 32'hc2cbbfa6} /* (23, 24, 3) {real, imag} */,
  {32'h44c3bc78, 32'h4355a464} /* (23, 24, 2) {real, imag} */,
  {32'hc57400dc, 32'hc402142f} /* (23, 24, 1) {real, imag} */,
  {32'hc579586c, 32'h00000000} /* (23, 24, 0) {real, imag} */,
  {32'hc54f85b2, 32'h43dbfe52} /* (23, 23, 31) {real, imag} */,
  {32'h44ab9ad8, 32'hc3079ce8} /* (23, 23, 30) {real, imag} */,
  {32'hc23dbe1c, 32'h422801c5} /* (23, 23, 29) {real, imag} */,
  {32'hc2af5581, 32'h42f89864} /* (23, 23, 28) {real, imag} */,
  {32'h43126ac2, 32'hc2a159ea} /* (23, 23, 27) {real, imag} */,
  {32'hc284dd79, 32'h41a259ae} /* (23, 23, 26) {real, imag} */,
  {32'hc1e19eb5, 32'h425c061a} /* (23, 23, 25) {real, imag} */,
  {32'hc235c3f2, 32'h42928923} /* (23, 23, 24) {real, imag} */,
  {32'hc231b02e, 32'h41891381} /* (23, 23, 23) {real, imag} */,
  {32'hc2280bc6, 32'h417ade8e} /* (23, 23, 22) {real, imag} */,
  {32'h42d07cc9, 32'hc255a092} /* (23, 23, 21) {real, imag} */,
  {32'hc06325b0, 32'h423bc5ef} /* (23, 23, 20) {real, imag} */,
  {32'h41997aec, 32'hc2d19f24} /* (23, 23, 19) {real, imag} */,
  {32'hc26b033e, 32'h420252c9} /* (23, 23, 18) {real, imag} */,
  {32'hc0705148, 32'h41c58f46} /* (23, 23, 17) {real, imag} */,
  {32'hc163c82a, 32'h00000000} /* (23, 23, 16) {real, imag} */,
  {32'hc0705148, 32'hc1c58f46} /* (23, 23, 15) {real, imag} */,
  {32'hc26b033e, 32'hc20252c9} /* (23, 23, 14) {real, imag} */,
  {32'h41997aec, 32'h42d19f24} /* (23, 23, 13) {real, imag} */,
  {32'hc06325b0, 32'hc23bc5ef} /* (23, 23, 12) {real, imag} */,
  {32'h42d07cc9, 32'h4255a092} /* (23, 23, 11) {real, imag} */,
  {32'hc2280bc6, 32'hc17ade8e} /* (23, 23, 10) {real, imag} */,
  {32'hc231b02e, 32'hc1891381} /* (23, 23, 9) {real, imag} */,
  {32'hc235c3f2, 32'hc2928923} /* (23, 23, 8) {real, imag} */,
  {32'hc1e19eb5, 32'hc25c061a} /* (23, 23, 7) {real, imag} */,
  {32'hc284dd79, 32'hc1a259ae} /* (23, 23, 6) {real, imag} */,
  {32'h43126ac2, 32'h42a159ea} /* (23, 23, 5) {real, imag} */,
  {32'hc2af5581, 32'hc2f89864} /* (23, 23, 4) {real, imag} */,
  {32'hc23dbe1c, 32'hc22801c5} /* (23, 23, 3) {real, imag} */,
  {32'h44ab9ad8, 32'h43079ce8} /* (23, 23, 2) {real, imag} */,
  {32'hc54f85b2, 32'hc3dbfe52} /* (23, 23, 1) {real, imag} */,
  {32'hc54422d6, 32'h00000000} /* (23, 23, 0) {real, imag} */,
  {32'hc512b5c2, 32'h436a84a1} /* (23, 22, 31) {real, imag} */,
  {32'h446c861f, 32'hc304baee} /* (23, 22, 30) {real, imag} */,
  {32'hc24f8e1a, 32'hc1bf0d6e} /* (23, 22, 29) {real, imag} */,
  {32'hc30c8ff3, 32'h43221bb6} /* (23, 22, 28) {real, imag} */,
  {32'h4354b0c5, 32'hc28feea9} /* (23, 22, 27) {real, imag} */,
  {32'hc2131dab, 32'h41dd3fc9} /* (23, 22, 26) {real, imag} */,
  {32'hc23cf9bc, 32'h4254d25c} /* (23, 22, 25) {real, imag} */,
  {32'h3fd39be0, 32'hc2a2cbca} /* (23, 22, 24) {real, imag} */,
  {32'hc29e025a, 32'h41c89ea5} /* (23, 22, 23) {real, imag} */,
  {32'h412c35dc, 32'hc1985c66} /* (23, 22, 22) {real, imag} */,
  {32'hc20914c4, 32'hc07eb3bc} /* (23, 22, 21) {real, imag} */,
  {32'h40e8f9f8, 32'hc13c0b60} /* (23, 22, 20) {real, imag} */,
  {32'hc20de986, 32'h3fd10fd0} /* (23, 22, 19) {real, imag} */,
  {32'h4283005e, 32'hc1cd53e2} /* (23, 22, 18) {real, imag} */,
  {32'hc1c7f47e, 32'hc18c0710} /* (23, 22, 17) {real, imag} */,
  {32'h41f23895, 32'h00000000} /* (23, 22, 16) {real, imag} */,
  {32'hc1c7f47e, 32'h418c0710} /* (23, 22, 15) {real, imag} */,
  {32'h4283005e, 32'h41cd53e2} /* (23, 22, 14) {real, imag} */,
  {32'hc20de986, 32'hbfd10fd0} /* (23, 22, 13) {real, imag} */,
  {32'h40e8f9f8, 32'h413c0b60} /* (23, 22, 12) {real, imag} */,
  {32'hc20914c4, 32'h407eb3bc} /* (23, 22, 11) {real, imag} */,
  {32'h412c35dc, 32'h41985c66} /* (23, 22, 10) {real, imag} */,
  {32'hc29e025a, 32'hc1c89ea5} /* (23, 22, 9) {real, imag} */,
  {32'h3fd39be0, 32'h42a2cbca} /* (23, 22, 8) {real, imag} */,
  {32'hc23cf9bc, 32'hc254d25c} /* (23, 22, 7) {real, imag} */,
  {32'hc2131dab, 32'hc1dd3fc9} /* (23, 22, 6) {real, imag} */,
  {32'h4354b0c5, 32'h428feea9} /* (23, 22, 5) {real, imag} */,
  {32'hc30c8ff3, 32'hc3221bb6} /* (23, 22, 4) {real, imag} */,
  {32'hc24f8e1a, 32'h41bf0d6e} /* (23, 22, 3) {real, imag} */,
  {32'h446c861f, 32'h4304baee} /* (23, 22, 2) {real, imag} */,
  {32'hc512b5c2, 32'hc36a84a1} /* (23, 22, 1) {real, imag} */,
  {32'hc5018be3, 32'h00000000} /* (23, 22, 0) {real, imag} */,
  {32'hc47c84a0, 32'h425e8188} /* (23, 21, 31) {real, imag} */,
  {32'h43acbe70, 32'hc3114a48} /* (23, 21, 30) {real, imag} */,
  {32'hc28c9901, 32'h42e97b94} /* (23, 21, 29) {real, imag} */,
  {32'h42388cff, 32'h42f373b8} /* (23, 21, 28) {real, imag} */,
  {32'h4328f298, 32'hc2a13113} /* (23, 21, 27) {real, imag} */,
  {32'hc295fc8f, 32'hc1e93855} /* (23, 21, 26) {real, imag} */,
  {32'h42e0c03a, 32'hc2d38f5c} /* (23, 21, 25) {real, imag} */,
  {32'hc316279e, 32'hc06f357c} /* (23, 21, 24) {real, imag} */,
  {32'hc28781e5, 32'hc246932e} /* (23, 21, 23) {real, imag} */,
  {32'hc209b5b6, 32'h42544839} /* (23, 21, 22) {real, imag} */,
  {32'h42c29761, 32'hc20425e6} /* (23, 21, 21) {real, imag} */,
  {32'hc23d7327, 32'hc19ee67b} /* (23, 21, 20) {real, imag} */,
  {32'hc2c731a1, 32'hc1aaf31c} /* (23, 21, 19) {real, imag} */,
  {32'h429d52ca, 32'hc0f43488} /* (23, 21, 18) {real, imag} */,
  {32'hc2557074, 32'h42272a58} /* (23, 21, 17) {real, imag} */,
  {32'hc03a8d00, 32'h00000000} /* (23, 21, 16) {real, imag} */,
  {32'hc2557074, 32'hc2272a58} /* (23, 21, 15) {real, imag} */,
  {32'h429d52ca, 32'h40f43488} /* (23, 21, 14) {real, imag} */,
  {32'hc2c731a1, 32'h41aaf31c} /* (23, 21, 13) {real, imag} */,
  {32'hc23d7327, 32'h419ee67b} /* (23, 21, 12) {real, imag} */,
  {32'h42c29761, 32'h420425e6} /* (23, 21, 11) {real, imag} */,
  {32'hc209b5b6, 32'hc2544839} /* (23, 21, 10) {real, imag} */,
  {32'hc28781e5, 32'h4246932e} /* (23, 21, 9) {real, imag} */,
  {32'hc316279e, 32'h406f357c} /* (23, 21, 8) {real, imag} */,
  {32'h42e0c03a, 32'h42d38f5c} /* (23, 21, 7) {real, imag} */,
  {32'hc295fc8f, 32'h41e93855} /* (23, 21, 6) {real, imag} */,
  {32'h4328f298, 32'h42a13113} /* (23, 21, 5) {real, imag} */,
  {32'h42388cff, 32'hc2f373b8} /* (23, 21, 4) {real, imag} */,
  {32'hc28c9901, 32'hc2e97b94} /* (23, 21, 3) {real, imag} */,
  {32'h43acbe70, 32'h43114a48} /* (23, 21, 2) {real, imag} */,
  {32'hc47c84a0, 32'hc25e8188} /* (23, 21, 1) {real, imag} */,
  {32'hc4876531, 32'h00000000} /* (23, 21, 0) {real, imag} */,
  {32'h44651645, 32'hc3204fa8} /* (23, 20, 31) {real, imag} */,
  {32'hc40a611c, 32'hc305eeff} /* (23, 20, 30) {real, imag} */,
  {32'hc13c41a0, 32'h432b06ee} /* (23, 20, 29) {real, imag} */,
  {32'h431d06e9, 32'hc3125ad9} /* (23, 20, 28) {real, imag} */,
  {32'hc1b12e40, 32'h4201dc90} /* (23, 20, 27) {real, imag} */,
  {32'hc3054b88, 32'hc2c0fc80} /* (23, 20, 26) {real, imag} */,
  {32'h425856a4, 32'hc2adb74a} /* (23, 20, 25) {real, imag} */,
  {32'hc32b4174, 32'h42391b56} /* (23, 20, 24) {real, imag} */,
  {32'h424e3659, 32'h4143497c} /* (23, 20, 23) {real, imag} */,
  {32'hc2721796, 32'hc18c020c} /* (23, 20, 22) {real, imag} */,
  {32'h430fa820, 32'h42ce54a7} /* (23, 20, 21) {real, imag} */,
  {32'hc26ebb44, 32'h40ca4a7c} /* (23, 20, 20) {real, imag} */,
  {32'hc26a2854, 32'h43029f96} /* (23, 20, 19) {real, imag} */,
  {32'h3e45fa00, 32'h426f83aa} /* (23, 20, 18) {real, imag} */,
  {32'hc1dcc77b, 32'hc0b3cd6c} /* (23, 20, 17) {real, imag} */,
  {32'hc1cc0d3c, 32'h00000000} /* (23, 20, 16) {real, imag} */,
  {32'hc1dcc77b, 32'h40b3cd6c} /* (23, 20, 15) {real, imag} */,
  {32'h3e45fa00, 32'hc26f83aa} /* (23, 20, 14) {real, imag} */,
  {32'hc26a2854, 32'hc3029f96} /* (23, 20, 13) {real, imag} */,
  {32'hc26ebb44, 32'hc0ca4a7c} /* (23, 20, 12) {real, imag} */,
  {32'h430fa820, 32'hc2ce54a7} /* (23, 20, 11) {real, imag} */,
  {32'hc2721796, 32'h418c020c} /* (23, 20, 10) {real, imag} */,
  {32'h424e3659, 32'hc143497c} /* (23, 20, 9) {real, imag} */,
  {32'hc32b4174, 32'hc2391b56} /* (23, 20, 8) {real, imag} */,
  {32'h425856a4, 32'h42adb74a} /* (23, 20, 7) {real, imag} */,
  {32'hc3054b88, 32'h42c0fc80} /* (23, 20, 6) {real, imag} */,
  {32'hc1b12e40, 32'hc201dc90} /* (23, 20, 5) {real, imag} */,
  {32'h431d06e9, 32'h43125ad9} /* (23, 20, 4) {real, imag} */,
  {32'hc13c41a0, 32'hc32b06ee} /* (23, 20, 3) {real, imag} */,
  {32'hc40a611c, 32'h4305eeff} /* (23, 20, 2) {real, imag} */,
  {32'h44651645, 32'h43204fa8} /* (23, 20, 1) {real, imag} */,
  {32'h43ef80ce, 32'h00000000} /* (23, 20, 0) {real, imag} */,
  {32'h4504e26f, 32'hc3a85f2d} /* (23, 19, 31) {real, imag} */,
  {32'hc446084e, 32'h43636225} /* (23, 19, 30) {real, imag} */,
  {32'hc1a62422, 32'h42d118ac} /* (23, 19, 29) {real, imag} */,
  {32'h4334c0a7, 32'hc393ab46} /* (23, 19, 28) {real, imag} */,
  {32'hc2e91676, 32'h41c68324} /* (23, 19, 27) {real, imag} */,
  {32'h413e65b8, 32'hc19cf768} /* (23, 19, 26) {real, imag} */,
  {32'h4262307f, 32'hc21b97dc} /* (23, 19, 25) {real, imag} */,
  {32'hc20c2a7a, 32'h4188fe91} /* (23, 19, 24) {real, imag} */,
  {32'hc2ab8f30, 32'h42b2c6aa} /* (23, 19, 23) {real, imag} */,
  {32'hc281fadd, 32'hc2017ac7} /* (23, 19, 22) {real, imag} */,
  {32'hc1bf95c0, 32'h41e391b2} /* (23, 19, 21) {real, imag} */,
  {32'hc2ef4c8b, 32'h4279a28e} /* (23, 19, 20) {real, imag} */,
  {32'h41a6d912, 32'hc1ca9216} /* (23, 19, 19) {real, imag} */,
  {32'h4081b1e8, 32'hc0bdaf78} /* (23, 19, 18) {real, imag} */,
  {32'h41d417bd, 32'h41a87aa1} /* (23, 19, 17) {real, imag} */,
  {32'hc10b3b36, 32'h00000000} /* (23, 19, 16) {real, imag} */,
  {32'h41d417bd, 32'hc1a87aa1} /* (23, 19, 15) {real, imag} */,
  {32'h4081b1e8, 32'h40bdaf78} /* (23, 19, 14) {real, imag} */,
  {32'h41a6d912, 32'h41ca9216} /* (23, 19, 13) {real, imag} */,
  {32'hc2ef4c8b, 32'hc279a28e} /* (23, 19, 12) {real, imag} */,
  {32'hc1bf95c0, 32'hc1e391b2} /* (23, 19, 11) {real, imag} */,
  {32'hc281fadd, 32'h42017ac7} /* (23, 19, 10) {real, imag} */,
  {32'hc2ab8f30, 32'hc2b2c6aa} /* (23, 19, 9) {real, imag} */,
  {32'hc20c2a7a, 32'hc188fe91} /* (23, 19, 8) {real, imag} */,
  {32'h4262307f, 32'h421b97dc} /* (23, 19, 7) {real, imag} */,
  {32'h413e65b8, 32'h419cf768} /* (23, 19, 6) {real, imag} */,
  {32'hc2e91676, 32'hc1c68324} /* (23, 19, 5) {real, imag} */,
  {32'h4334c0a7, 32'h4393ab46} /* (23, 19, 4) {real, imag} */,
  {32'hc1a62422, 32'hc2d118ac} /* (23, 19, 3) {real, imag} */,
  {32'hc446084e, 32'hc3636225} /* (23, 19, 2) {real, imag} */,
  {32'h4504e26f, 32'h43a85f2d} /* (23, 19, 1) {real, imag} */,
  {32'h44af93c8, 32'h00000000} /* (23, 19, 0) {real, imag} */,
  {32'h453a755a, 32'hc38aeb90} /* (23, 18, 31) {real, imag} */,
  {32'hc485029c, 32'h4383646e} /* (23, 18, 30) {real, imag} */,
  {32'h40debb10, 32'h41b1a6f9} /* (23, 18, 29) {real, imag} */,
  {32'h439fca81, 32'hc3772bf6} /* (23, 18, 28) {real, imag} */,
  {32'hc39e73d8, 32'h4286bbb2} /* (23, 18, 27) {real, imag} */,
  {32'h42956017, 32'h428ae5a3} /* (23, 18, 26) {real, imag} */,
  {32'hc23cba30, 32'h41def434} /* (23, 18, 25) {real, imag} */,
  {32'h40e91978, 32'h4319c1db} /* (23, 18, 24) {real, imag} */,
  {32'hc0f12f1f, 32'h419dd4fb} /* (23, 18, 23) {real, imag} */,
  {32'hc20db31c, 32'h42d25e9e} /* (23, 18, 22) {real, imag} */,
  {32'h40745818, 32'h42c4e476} /* (23, 18, 21) {real, imag} */,
  {32'hc165d736, 32'hc1e0aa8a} /* (23, 18, 20) {real, imag} */,
  {32'h42687e9c, 32'h41515586} /* (23, 18, 19) {real, imag} */,
  {32'hc1aa285d, 32'h41dfcd9b} /* (23, 18, 18) {real, imag} */,
  {32'hc1ed5694, 32'hc251e129} /* (23, 18, 17) {real, imag} */,
  {32'hc1dc6df0, 32'h00000000} /* (23, 18, 16) {real, imag} */,
  {32'hc1ed5694, 32'h4251e129} /* (23, 18, 15) {real, imag} */,
  {32'hc1aa285d, 32'hc1dfcd9b} /* (23, 18, 14) {real, imag} */,
  {32'h42687e9c, 32'hc1515586} /* (23, 18, 13) {real, imag} */,
  {32'hc165d736, 32'h41e0aa8a} /* (23, 18, 12) {real, imag} */,
  {32'h40745818, 32'hc2c4e476} /* (23, 18, 11) {real, imag} */,
  {32'hc20db31c, 32'hc2d25e9e} /* (23, 18, 10) {real, imag} */,
  {32'hc0f12f1f, 32'hc19dd4fb} /* (23, 18, 9) {real, imag} */,
  {32'h40e91978, 32'hc319c1db} /* (23, 18, 8) {real, imag} */,
  {32'hc23cba30, 32'hc1def434} /* (23, 18, 7) {real, imag} */,
  {32'h42956017, 32'hc28ae5a3} /* (23, 18, 6) {real, imag} */,
  {32'hc39e73d8, 32'hc286bbb2} /* (23, 18, 5) {real, imag} */,
  {32'h439fca81, 32'h43772bf6} /* (23, 18, 4) {real, imag} */,
  {32'h40debb10, 32'hc1b1a6f9} /* (23, 18, 3) {real, imag} */,
  {32'hc485029c, 32'hc383646e} /* (23, 18, 2) {real, imag} */,
  {32'h453a755a, 32'h438aeb90} /* (23, 18, 1) {real, imag} */,
  {32'h44f075c4, 32'h00000000} /* (23, 18, 0) {real, imag} */,
  {32'h455eef41, 32'hc3b4a511} /* (23, 17, 31) {real, imag} */,
  {32'hc49534c8, 32'h439be5d7} /* (23, 17, 30) {real, imag} */,
  {32'h4216ce4e, 32'hc12499c8} /* (23, 17, 29) {real, imag} */,
  {32'h43bf64e7, 32'hc383b61b} /* (23, 17, 28) {real, imag} */,
  {32'hc33b185a, 32'h42b8cb2f} /* (23, 17, 27) {real, imag} */,
  {32'hc289bcd7, 32'h42254944} /* (23, 17, 26) {real, imag} */,
  {32'h4222e8d4, 32'hc1ff5356} /* (23, 17, 25) {real, imag} */,
  {32'h4238b8a7, 32'h42d2e44c} /* (23, 17, 24) {real, imag} */,
  {32'hc1df9222, 32'hc21999f0} /* (23, 17, 23) {real, imag} */,
  {32'h41cdcefe, 32'hc309e442} /* (23, 17, 22) {real, imag} */,
  {32'hc2979034, 32'h41387891} /* (23, 17, 21) {real, imag} */,
  {32'h3f2a52c0, 32'h4191f8bb} /* (23, 17, 20) {real, imag} */,
  {32'hc2c0142a, 32'h422694ae} /* (23, 17, 19) {real, imag} */,
  {32'hc194509b, 32'h42a1e943} /* (23, 17, 18) {real, imag} */,
  {32'h41a48631, 32'hc0c23ab4} /* (23, 17, 17) {real, imag} */,
  {32'hc16607fa, 32'h00000000} /* (23, 17, 16) {real, imag} */,
  {32'h41a48631, 32'h40c23ab4} /* (23, 17, 15) {real, imag} */,
  {32'hc194509b, 32'hc2a1e943} /* (23, 17, 14) {real, imag} */,
  {32'hc2c0142a, 32'hc22694ae} /* (23, 17, 13) {real, imag} */,
  {32'h3f2a52c0, 32'hc191f8bb} /* (23, 17, 12) {real, imag} */,
  {32'hc2979034, 32'hc1387891} /* (23, 17, 11) {real, imag} */,
  {32'h41cdcefe, 32'h4309e442} /* (23, 17, 10) {real, imag} */,
  {32'hc1df9222, 32'h421999f0} /* (23, 17, 9) {real, imag} */,
  {32'h4238b8a7, 32'hc2d2e44c} /* (23, 17, 8) {real, imag} */,
  {32'h4222e8d4, 32'h41ff5356} /* (23, 17, 7) {real, imag} */,
  {32'hc289bcd7, 32'hc2254944} /* (23, 17, 6) {real, imag} */,
  {32'hc33b185a, 32'hc2b8cb2f} /* (23, 17, 5) {real, imag} */,
  {32'h43bf64e7, 32'h4383b61b} /* (23, 17, 4) {real, imag} */,
  {32'h4216ce4e, 32'h412499c8} /* (23, 17, 3) {real, imag} */,
  {32'hc49534c8, 32'hc39be5d7} /* (23, 17, 2) {real, imag} */,
  {32'h455eef41, 32'h43b4a511} /* (23, 17, 1) {real, imag} */,
  {32'h4505a853, 32'h00000000} /* (23, 17, 0) {real, imag} */,
  {32'h4568c5ee, 32'hc3cbf708} /* (23, 16, 31) {real, imag} */,
  {32'hc4a0c1dd, 32'h43a30785} /* (23, 16, 30) {real, imag} */,
  {32'h41cc402a, 32'h42d67ffc} /* (23, 16, 29) {real, imag} */,
  {32'h43a548a6, 32'hc30d8802} /* (23, 16, 28) {real, imag} */,
  {32'hc38288d2, 32'h42a30f6d} /* (23, 16, 27) {real, imag} */,
  {32'hc30a9bd1, 32'hc0834470} /* (23, 16, 26) {real, imag} */,
  {32'h42d1c41a, 32'hc0894d78} /* (23, 16, 25) {real, imag} */,
  {32'hc29b74a6, 32'h42c32716} /* (23, 16, 24) {real, imag} */,
  {32'hc285db8c, 32'h42c31e25} /* (23, 16, 23) {real, imag} */,
  {32'hc0c31545, 32'hc192d176} /* (23, 16, 22) {real, imag} */,
  {32'hc25e0010, 32'h41577865} /* (23, 16, 21) {real, imag} */,
  {32'hc212de2b, 32'h41835090} /* (23, 16, 20) {real, imag} */,
  {32'h41856ba4, 32'hc2861b2e} /* (23, 16, 19) {real, imag} */,
  {32'h42516b20, 32'hc2a38b0c} /* (23, 16, 18) {real, imag} */,
  {32'h4171304a, 32'hc1202802} /* (23, 16, 17) {real, imag} */,
  {32'hc2c573be, 32'h00000000} /* (23, 16, 16) {real, imag} */,
  {32'h4171304a, 32'h41202802} /* (23, 16, 15) {real, imag} */,
  {32'h42516b20, 32'h42a38b0c} /* (23, 16, 14) {real, imag} */,
  {32'h41856ba4, 32'h42861b2e} /* (23, 16, 13) {real, imag} */,
  {32'hc212de2b, 32'hc1835090} /* (23, 16, 12) {real, imag} */,
  {32'hc25e0010, 32'hc1577865} /* (23, 16, 11) {real, imag} */,
  {32'hc0c31545, 32'h4192d176} /* (23, 16, 10) {real, imag} */,
  {32'hc285db8c, 32'hc2c31e25} /* (23, 16, 9) {real, imag} */,
  {32'hc29b74a6, 32'hc2c32716} /* (23, 16, 8) {real, imag} */,
  {32'h42d1c41a, 32'h40894d78} /* (23, 16, 7) {real, imag} */,
  {32'hc30a9bd1, 32'h40834470} /* (23, 16, 6) {real, imag} */,
  {32'hc38288d2, 32'hc2a30f6d} /* (23, 16, 5) {real, imag} */,
  {32'h43a548a6, 32'h430d8802} /* (23, 16, 4) {real, imag} */,
  {32'h41cc402a, 32'hc2d67ffc} /* (23, 16, 3) {real, imag} */,
  {32'hc4a0c1dd, 32'hc3a30785} /* (23, 16, 2) {real, imag} */,
  {32'h4568c5ee, 32'h43cbf708} /* (23, 16, 1) {real, imag} */,
  {32'h451d55d4, 32'h00000000} /* (23, 16, 0) {real, imag} */,
  {32'h456cff65, 32'hc3977057} /* (23, 15, 31) {real, imag} */,
  {32'hc4a2f2c0, 32'h435407aa} /* (23, 15, 30) {real, imag} */,
  {32'hc32d85fe, 32'h42e1fa41} /* (23, 15, 29) {real, imag} */,
  {32'h438c12b1, 32'hc2c3f174} /* (23, 15, 28) {real, imag} */,
  {32'hc372dc1a, 32'h42e1f2f5} /* (23, 15, 27) {real, imag} */,
  {32'hc1137ca8, 32'hc21a7ba8} /* (23, 15, 26) {real, imag} */,
  {32'h42aab047, 32'hc1770f9c} /* (23, 15, 25) {real, imag} */,
  {32'hc31a1afa, 32'hc2b76228} /* (23, 15, 24) {real, imag} */,
  {32'h412155f4, 32'h42bc7f02} /* (23, 15, 23) {real, imag} */,
  {32'h40887aa2, 32'h42782916} /* (23, 15, 22) {real, imag} */,
  {32'h423dbf5c, 32'hc1b5e8ee} /* (23, 15, 21) {real, imag} */,
  {32'h42d59b6c, 32'h422de9a4} /* (23, 15, 20) {real, imag} */,
  {32'hc1fe3850, 32'hc2ea3941} /* (23, 15, 19) {real, imag} */,
  {32'h3d8e0100, 32'h41dc77c0} /* (23, 15, 18) {real, imag} */,
  {32'h41c6bea9, 32'hc2448a00} /* (23, 15, 17) {real, imag} */,
  {32'hc28929a9, 32'h00000000} /* (23, 15, 16) {real, imag} */,
  {32'h41c6bea9, 32'h42448a00} /* (23, 15, 15) {real, imag} */,
  {32'h3d8e0100, 32'hc1dc77c0} /* (23, 15, 14) {real, imag} */,
  {32'hc1fe3850, 32'h42ea3941} /* (23, 15, 13) {real, imag} */,
  {32'h42d59b6c, 32'hc22de9a4} /* (23, 15, 12) {real, imag} */,
  {32'h423dbf5c, 32'h41b5e8ee} /* (23, 15, 11) {real, imag} */,
  {32'h40887aa2, 32'hc2782916} /* (23, 15, 10) {real, imag} */,
  {32'h412155f4, 32'hc2bc7f02} /* (23, 15, 9) {real, imag} */,
  {32'hc31a1afa, 32'h42b76228} /* (23, 15, 8) {real, imag} */,
  {32'h42aab047, 32'h41770f9c} /* (23, 15, 7) {real, imag} */,
  {32'hc1137ca8, 32'h421a7ba8} /* (23, 15, 6) {real, imag} */,
  {32'hc372dc1a, 32'hc2e1f2f5} /* (23, 15, 5) {real, imag} */,
  {32'h438c12b1, 32'h42c3f174} /* (23, 15, 4) {real, imag} */,
  {32'hc32d85fe, 32'hc2e1fa41} /* (23, 15, 3) {real, imag} */,
  {32'hc4a2f2c0, 32'hc35407aa} /* (23, 15, 2) {real, imag} */,
  {32'h456cff65, 32'h43977057} /* (23, 15, 1) {real, imag} */,
  {32'h45205b67, 32'h00000000} /* (23, 15, 0) {real, imag} */,
  {32'h4555db62, 32'hc2db9320} /* (23, 14, 31) {real, imag} */,
  {32'hc4ab1dd8, 32'h43629c5f} /* (23, 14, 30) {real, imag} */,
  {32'hc2afe72d, 32'h4237febc} /* (23, 14, 29) {real, imag} */,
  {32'h43b2d9d7, 32'hc35834be} /* (23, 14, 28) {real, imag} */,
  {32'hc3756034, 32'h427dd9d3} /* (23, 14, 27) {real, imag} */,
  {32'hc2d2bfed, 32'h401ed460} /* (23, 14, 26) {real, imag} */,
  {32'h42f1d47e, 32'hc23114da} /* (23, 14, 25) {real, imag} */,
  {32'h42c390a8, 32'hc22825c5} /* (23, 14, 24) {real, imag} */,
  {32'h41457e68, 32'hc1314e62} /* (23, 14, 23) {real, imag} */,
  {32'h4067b1f8, 32'h42210ef7} /* (23, 14, 22) {real, imag} */,
  {32'hc1895fdd, 32'h42a2021e} /* (23, 14, 21) {real, imag} */,
  {32'h420e2170, 32'hc264afc7} /* (23, 14, 20) {real, imag} */,
  {32'h4209c000, 32'h423c0f12} /* (23, 14, 19) {real, imag} */,
  {32'hc1ff85ff, 32'h422e5ca2} /* (23, 14, 18) {real, imag} */,
  {32'h41278d9b, 32'h41ddb7d2} /* (23, 14, 17) {real, imag} */,
  {32'h42082dcb, 32'h00000000} /* (23, 14, 16) {real, imag} */,
  {32'h41278d9b, 32'hc1ddb7d2} /* (23, 14, 15) {real, imag} */,
  {32'hc1ff85ff, 32'hc22e5ca2} /* (23, 14, 14) {real, imag} */,
  {32'h4209c000, 32'hc23c0f12} /* (23, 14, 13) {real, imag} */,
  {32'h420e2170, 32'h4264afc7} /* (23, 14, 12) {real, imag} */,
  {32'hc1895fdd, 32'hc2a2021e} /* (23, 14, 11) {real, imag} */,
  {32'h4067b1f8, 32'hc2210ef7} /* (23, 14, 10) {real, imag} */,
  {32'h41457e68, 32'h41314e62} /* (23, 14, 9) {real, imag} */,
  {32'h42c390a8, 32'h422825c5} /* (23, 14, 8) {real, imag} */,
  {32'h42f1d47e, 32'h423114da} /* (23, 14, 7) {real, imag} */,
  {32'hc2d2bfed, 32'hc01ed460} /* (23, 14, 6) {real, imag} */,
  {32'hc3756034, 32'hc27dd9d3} /* (23, 14, 5) {real, imag} */,
  {32'h43b2d9d7, 32'h435834be} /* (23, 14, 4) {real, imag} */,
  {32'hc2afe72d, 32'hc237febc} /* (23, 14, 3) {real, imag} */,
  {32'hc4ab1dd8, 32'hc3629c5f} /* (23, 14, 2) {real, imag} */,
  {32'h4555db62, 32'h42db9320} /* (23, 14, 1) {real, imag} */,
  {32'h4522e7e0, 32'h00000000} /* (23, 14, 0) {real, imag} */,
  {32'h45351305, 32'hc258ea98} /* (23, 13, 31) {real, imag} */,
  {32'hc4ad1131, 32'h43231c1f} /* (23, 13, 30) {real, imag} */,
  {32'hc2ae87e8, 32'hc11f4f90} /* (23, 13, 29) {real, imag} */,
  {32'h43a13e0c, 32'hc398083c} /* (23, 13, 28) {real, imag} */,
  {32'hc391c26a, 32'h4302a688} /* (23, 13, 27) {real, imag} */,
  {32'h42a787e3, 32'h41a2a9a4} /* (23, 13, 26) {real, imag} */,
  {32'h433569e3, 32'h4250d1d2} /* (23, 13, 25) {real, imag} */,
  {32'hc005e9a0, 32'hc1536cf2} /* (23, 13, 24) {real, imag} */,
  {32'h42a7fdac, 32'h410a7d60} /* (23, 13, 23) {real, imag} */,
  {32'h40c835bc, 32'h40b486f8} /* (23, 13, 22) {real, imag} */,
  {32'h42882d14, 32'h42b50654} /* (23, 13, 21) {real, imag} */,
  {32'h40bb4c50, 32'h4187b8f4} /* (23, 13, 20) {real, imag} */,
  {32'hc293d4cc, 32'hc1e11a60} /* (23, 13, 19) {real, imag} */,
  {32'h4219298d, 32'hc222c123} /* (23, 13, 18) {real, imag} */,
  {32'hc2895245, 32'h417e8f42} /* (23, 13, 17) {real, imag} */,
  {32'hc2434c56, 32'h00000000} /* (23, 13, 16) {real, imag} */,
  {32'hc2895245, 32'hc17e8f42} /* (23, 13, 15) {real, imag} */,
  {32'h4219298d, 32'h4222c123} /* (23, 13, 14) {real, imag} */,
  {32'hc293d4cc, 32'h41e11a60} /* (23, 13, 13) {real, imag} */,
  {32'h40bb4c50, 32'hc187b8f4} /* (23, 13, 12) {real, imag} */,
  {32'h42882d14, 32'hc2b50654} /* (23, 13, 11) {real, imag} */,
  {32'h40c835bc, 32'hc0b486f8} /* (23, 13, 10) {real, imag} */,
  {32'h42a7fdac, 32'hc10a7d60} /* (23, 13, 9) {real, imag} */,
  {32'hc005e9a0, 32'h41536cf2} /* (23, 13, 8) {real, imag} */,
  {32'h433569e3, 32'hc250d1d2} /* (23, 13, 7) {real, imag} */,
  {32'h42a787e3, 32'hc1a2a9a4} /* (23, 13, 6) {real, imag} */,
  {32'hc391c26a, 32'hc302a688} /* (23, 13, 5) {real, imag} */,
  {32'h43a13e0c, 32'h4398083c} /* (23, 13, 4) {real, imag} */,
  {32'hc2ae87e8, 32'h411f4f90} /* (23, 13, 3) {real, imag} */,
  {32'hc4ad1131, 32'hc3231c1f} /* (23, 13, 2) {real, imag} */,
  {32'h45351305, 32'h4258ea98} /* (23, 13, 1) {real, imag} */,
  {32'h4508f8be, 32'h00000000} /* (23, 13, 0) {real, imag} */,
  {32'h45147b31, 32'h4334fe98} /* (23, 12, 31) {real, imag} */,
  {32'hc4928008, 32'h42d2b5d2} /* (23, 12, 30) {real, imag} */,
  {32'hc2842e50, 32'h411fd7e0} /* (23, 12, 29) {real, imag} */,
  {32'h438712dc, 32'hc3737d13} /* (23, 12, 28) {real, imag} */,
  {32'hc349c80e, 32'h4398aea4} /* (23, 12, 27) {real, imag} */,
  {32'h416fc3a4, 32'hc29a73a0} /* (23, 12, 26) {real, imag} */,
  {32'h42ec5088, 32'hc1b4305c} /* (23, 12, 25) {real, imag} */,
  {32'hc3053afc, 32'h41aae8f0} /* (23, 12, 24) {real, imag} */,
  {32'hc20bd3f9, 32'h42933e2e} /* (23, 12, 23) {real, imag} */,
  {32'h4226b924, 32'hc28bf754} /* (23, 12, 22) {real, imag} */,
  {32'hc1d5b642, 32'hc20fa8a2} /* (23, 12, 21) {real, imag} */,
  {32'hc0947760, 32'hc1d34e53} /* (23, 12, 20) {real, imag} */,
  {32'hc01f2dd8, 32'hc21a4232} /* (23, 12, 19) {real, imag} */,
  {32'hc2168159, 32'h42b133f3} /* (23, 12, 18) {real, imag} */,
  {32'hc1d4c067, 32'h4202f98e} /* (23, 12, 17) {real, imag} */,
  {32'h42c64e15, 32'h00000000} /* (23, 12, 16) {real, imag} */,
  {32'hc1d4c067, 32'hc202f98e} /* (23, 12, 15) {real, imag} */,
  {32'hc2168159, 32'hc2b133f3} /* (23, 12, 14) {real, imag} */,
  {32'hc01f2dd8, 32'h421a4232} /* (23, 12, 13) {real, imag} */,
  {32'hc0947760, 32'h41d34e53} /* (23, 12, 12) {real, imag} */,
  {32'hc1d5b642, 32'h420fa8a2} /* (23, 12, 11) {real, imag} */,
  {32'h4226b924, 32'h428bf754} /* (23, 12, 10) {real, imag} */,
  {32'hc20bd3f9, 32'hc2933e2e} /* (23, 12, 9) {real, imag} */,
  {32'hc3053afc, 32'hc1aae8f0} /* (23, 12, 8) {real, imag} */,
  {32'h42ec5088, 32'h41b4305c} /* (23, 12, 7) {real, imag} */,
  {32'h416fc3a4, 32'h429a73a0} /* (23, 12, 6) {real, imag} */,
  {32'hc349c80e, 32'hc398aea4} /* (23, 12, 5) {real, imag} */,
  {32'h438712dc, 32'h43737d13} /* (23, 12, 4) {real, imag} */,
  {32'hc2842e50, 32'hc11fd7e0} /* (23, 12, 3) {real, imag} */,
  {32'hc4928008, 32'hc2d2b5d2} /* (23, 12, 2) {real, imag} */,
  {32'h45147b31, 32'hc334fe98} /* (23, 12, 1) {real, imag} */,
  {32'h44bd5ca4, 32'h00000000} /* (23, 12, 0) {real, imag} */,
  {32'h4495d2fc, 32'h4359ea6e} /* (23, 11, 31) {real, imag} */,
  {32'hc438e32a, 32'hc2b4b46f} /* (23, 11, 30) {real, imag} */,
  {32'hc33a60c0, 32'hc1797c24} /* (23, 11, 29) {real, imag} */,
  {32'h432a69bc, 32'hc27d1f68} /* (23, 11, 28) {real, imag} */,
  {32'hc338138c, 32'h42f3a763} /* (23, 11, 27) {real, imag} */,
  {32'hc26c0231, 32'h41ab3da3} /* (23, 11, 26) {real, imag} */,
  {32'h4295a0a8, 32'hc03f1f00} /* (23, 11, 25) {real, imag} */,
  {32'hc299af60, 32'h40de940a} /* (23, 11, 24) {real, imag} */,
  {32'h41f6e655, 32'hc28ed31f} /* (23, 11, 23) {real, imag} */,
  {32'hc140605a, 32'hc1eb3b8e} /* (23, 11, 22) {real, imag} */,
  {32'hc2350716, 32'h425f210a} /* (23, 11, 21) {real, imag} */,
  {32'hc242bc65, 32'hc030ac08} /* (23, 11, 20) {real, imag} */,
  {32'hc26f1ba2, 32'h4206d379} /* (23, 11, 19) {real, imag} */,
  {32'h41d482e4, 32'hc2875c1e} /* (23, 11, 18) {real, imag} */,
  {32'h41afc5c0, 32'h4146e1ac} /* (23, 11, 17) {real, imag} */,
  {32'h42b7f5b3, 32'h00000000} /* (23, 11, 16) {real, imag} */,
  {32'h41afc5c0, 32'hc146e1ac} /* (23, 11, 15) {real, imag} */,
  {32'h41d482e4, 32'h42875c1e} /* (23, 11, 14) {real, imag} */,
  {32'hc26f1ba2, 32'hc206d379} /* (23, 11, 13) {real, imag} */,
  {32'hc242bc65, 32'h4030ac08} /* (23, 11, 12) {real, imag} */,
  {32'hc2350716, 32'hc25f210a} /* (23, 11, 11) {real, imag} */,
  {32'hc140605a, 32'h41eb3b8e} /* (23, 11, 10) {real, imag} */,
  {32'h41f6e655, 32'h428ed31f} /* (23, 11, 9) {real, imag} */,
  {32'hc299af60, 32'hc0de940a} /* (23, 11, 8) {real, imag} */,
  {32'h4295a0a8, 32'h403f1f00} /* (23, 11, 7) {real, imag} */,
  {32'hc26c0231, 32'hc1ab3da3} /* (23, 11, 6) {real, imag} */,
  {32'hc338138c, 32'hc2f3a763} /* (23, 11, 5) {real, imag} */,
  {32'h432a69bc, 32'h427d1f68} /* (23, 11, 4) {real, imag} */,
  {32'hc33a60c0, 32'h41797c24} /* (23, 11, 3) {real, imag} */,
  {32'hc438e32a, 32'h42b4b46f} /* (23, 11, 2) {real, imag} */,
  {32'h4495d2fc, 32'hc359ea6e} /* (23, 11, 1) {real, imag} */,
  {32'h4408ef3a, 32'h00000000} /* (23, 11, 0) {real, imag} */,
  {32'hc424b28f, 32'h4415887a} /* (23, 10, 31) {real, imag} */,
  {32'h4080fa80, 32'hc3aff770} /* (23, 10, 30) {real, imag} */,
  {32'hc32e0572, 32'hc25c8e4b} /* (23, 10, 29) {real, imag} */,
  {32'h434e6633, 32'h42b3b628} /* (23, 10, 28) {real, imag} */,
  {32'h4309e1d7, 32'hc29a4a7b} /* (23, 10, 27) {real, imag} */,
  {32'hc09e4086, 32'hc13bfdde} /* (23, 10, 26) {real, imag} */,
  {32'hc29d417a, 32'h41e02c60} /* (23, 10, 25) {real, imag} */,
  {32'h42ced292, 32'h430e4823} /* (23, 10, 24) {real, imag} */,
  {32'h42236099, 32'h420faa44} /* (23, 10, 23) {real, imag} */,
  {32'hc2a2a876, 32'hc2a0bc42} /* (23, 10, 22) {real, imag} */,
  {32'hc26cfc7e, 32'hc0ac7abe} /* (23, 10, 21) {real, imag} */,
  {32'h423646c0, 32'hc14c46a4} /* (23, 10, 20) {real, imag} */,
  {32'h4214af44, 32'hc259fff6} /* (23, 10, 19) {real, imag} */,
  {32'h41ce8a88, 32'hc21d99a7} /* (23, 10, 18) {real, imag} */,
  {32'h41ded882, 32'h42a55c2e} /* (23, 10, 17) {real, imag} */,
  {32'h4294b030, 32'h00000000} /* (23, 10, 16) {real, imag} */,
  {32'h41ded882, 32'hc2a55c2e} /* (23, 10, 15) {real, imag} */,
  {32'h41ce8a88, 32'h421d99a7} /* (23, 10, 14) {real, imag} */,
  {32'h4214af44, 32'h4259fff6} /* (23, 10, 13) {real, imag} */,
  {32'h423646c0, 32'h414c46a4} /* (23, 10, 12) {real, imag} */,
  {32'hc26cfc7e, 32'h40ac7abe} /* (23, 10, 11) {real, imag} */,
  {32'hc2a2a876, 32'h42a0bc42} /* (23, 10, 10) {real, imag} */,
  {32'h42236099, 32'hc20faa44} /* (23, 10, 9) {real, imag} */,
  {32'h42ced292, 32'hc30e4823} /* (23, 10, 8) {real, imag} */,
  {32'hc29d417a, 32'hc1e02c60} /* (23, 10, 7) {real, imag} */,
  {32'hc09e4086, 32'h413bfdde} /* (23, 10, 6) {real, imag} */,
  {32'h4309e1d7, 32'h429a4a7b} /* (23, 10, 5) {real, imag} */,
  {32'h434e6633, 32'hc2b3b628} /* (23, 10, 4) {real, imag} */,
  {32'hc32e0572, 32'h425c8e4b} /* (23, 10, 3) {real, imag} */,
  {32'h4080fa80, 32'h43aff770} /* (23, 10, 2) {real, imag} */,
  {32'hc424b28f, 32'hc415887a} /* (23, 10, 1) {real, imag} */,
  {32'hc4625ccf, 32'h00000000} /* (23, 10, 0) {real, imag} */,
  {32'hc4f6a76c, 32'h4484d124} /* (23, 9, 31) {real, imag} */,
  {32'h442e194f, 32'hc396a720} /* (23, 9, 30) {real, imag} */,
  {32'hc29d620e, 32'h42cbbb5c} /* (23, 9, 29) {real, imag} */,
  {32'hc18bc84c, 32'h42896fda} /* (23, 9, 28) {real, imag} */,
  {32'h4369171c, 32'hc2624dc8} /* (23, 9, 27) {real, imag} */,
  {32'h424c3a56, 32'hc082ac46} /* (23, 9, 26) {real, imag} */,
  {32'h42042977, 32'hc1c935ac} /* (23, 9, 25) {real, imag} */,
  {32'h42a55689, 32'hc2526ea6} /* (23, 9, 24) {real, imag} */,
  {32'h41d45627, 32'h41eccbcf} /* (23, 9, 23) {real, imag} */,
  {32'hc1803ebe, 32'h423f9ce4} /* (23, 9, 22) {real, imag} */,
  {32'h429a8f13, 32'h41a898f8} /* (23, 9, 21) {real, imag} */,
  {32'hc29dd556, 32'h422c81b9} /* (23, 9, 20) {real, imag} */,
  {32'hc24a722e, 32'hc10b63f4} /* (23, 9, 19) {real, imag} */,
  {32'hc18900bd, 32'hc08d71aa} /* (23, 9, 18) {real, imag} */,
  {32'h421fe26a, 32'h41d2ae6e} /* (23, 9, 17) {real, imag} */,
  {32'hc2756e60, 32'h00000000} /* (23, 9, 16) {real, imag} */,
  {32'h421fe26a, 32'hc1d2ae6e} /* (23, 9, 15) {real, imag} */,
  {32'hc18900bd, 32'h408d71aa} /* (23, 9, 14) {real, imag} */,
  {32'hc24a722e, 32'h410b63f4} /* (23, 9, 13) {real, imag} */,
  {32'hc29dd556, 32'hc22c81b9} /* (23, 9, 12) {real, imag} */,
  {32'h429a8f13, 32'hc1a898f8} /* (23, 9, 11) {real, imag} */,
  {32'hc1803ebe, 32'hc23f9ce4} /* (23, 9, 10) {real, imag} */,
  {32'h41d45627, 32'hc1eccbcf} /* (23, 9, 9) {real, imag} */,
  {32'h42a55689, 32'h42526ea6} /* (23, 9, 8) {real, imag} */,
  {32'h42042977, 32'h41c935ac} /* (23, 9, 7) {real, imag} */,
  {32'h424c3a56, 32'h4082ac46} /* (23, 9, 6) {real, imag} */,
  {32'h4369171c, 32'h42624dc8} /* (23, 9, 5) {real, imag} */,
  {32'hc18bc84c, 32'hc2896fda} /* (23, 9, 4) {real, imag} */,
  {32'hc29d620e, 32'hc2cbbb5c} /* (23, 9, 3) {real, imag} */,
  {32'h442e194f, 32'h4396a720} /* (23, 9, 2) {real, imag} */,
  {32'hc4f6a76c, 32'hc484d124} /* (23, 9, 1) {real, imag} */,
  {32'hc50b7d1a, 32'h00000000} /* (23, 9, 0) {real, imag} */,
  {32'hc530b814, 32'h44b8ab3e} /* (23, 8, 31) {real, imag} */,
  {32'h446316c7, 32'hc3e5fbc0} /* (23, 8, 30) {real, imag} */,
  {32'h4318f415, 32'h42b5d76a} /* (23, 8, 29) {real, imag} */,
  {32'hc30eedc1, 32'h42b2339f} /* (23, 8, 28) {real, imag} */,
  {32'h433c80c4, 32'hc2fe296b} /* (23, 8, 27) {real, imag} */,
  {32'h42fa7be8, 32'hc1a6c0f6} /* (23, 8, 26) {real, imag} */,
  {32'hc2885378, 32'h429fe3e0} /* (23, 8, 25) {real, imag} */,
  {32'h427ade62, 32'h41500b94} /* (23, 8, 24) {real, imag} */,
  {32'hc2e21a72, 32'h42877aa7} /* (23, 8, 23) {real, imag} */,
  {32'h42034a9d, 32'hc3044ffd} /* (23, 8, 22) {real, imag} */,
  {32'h423fd98b, 32'h4215ef3a} /* (23, 8, 21) {real, imag} */,
  {32'hc324ce81, 32'hc26ccff8} /* (23, 8, 20) {real, imag} */,
  {32'h420c7552, 32'h424483bd} /* (23, 8, 19) {real, imag} */,
  {32'h4124a210, 32'hc2451633} /* (23, 8, 18) {real, imag} */,
  {32'h41a92d00, 32'hc23a8a0a} /* (23, 8, 17) {real, imag} */,
  {32'h420b68c1, 32'h00000000} /* (23, 8, 16) {real, imag} */,
  {32'h41a92d00, 32'h423a8a0a} /* (23, 8, 15) {real, imag} */,
  {32'h4124a210, 32'h42451633} /* (23, 8, 14) {real, imag} */,
  {32'h420c7552, 32'hc24483bd} /* (23, 8, 13) {real, imag} */,
  {32'hc324ce81, 32'h426ccff8} /* (23, 8, 12) {real, imag} */,
  {32'h423fd98b, 32'hc215ef3a} /* (23, 8, 11) {real, imag} */,
  {32'h42034a9d, 32'h43044ffd} /* (23, 8, 10) {real, imag} */,
  {32'hc2e21a72, 32'hc2877aa7} /* (23, 8, 9) {real, imag} */,
  {32'h427ade62, 32'hc1500b94} /* (23, 8, 8) {real, imag} */,
  {32'hc2885378, 32'hc29fe3e0} /* (23, 8, 7) {real, imag} */,
  {32'h42fa7be8, 32'h41a6c0f6} /* (23, 8, 6) {real, imag} */,
  {32'h433c80c4, 32'h42fe296b} /* (23, 8, 5) {real, imag} */,
  {32'hc30eedc1, 32'hc2b2339f} /* (23, 8, 4) {real, imag} */,
  {32'h4318f415, 32'hc2b5d76a} /* (23, 8, 3) {real, imag} */,
  {32'h446316c7, 32'h43e5fbc0} /* (23, 8, 2) {real, imag} */,
  {32'hc530b814, 32'hc4b8ab3e} /* (23, 8, 1) {real, imag} */,
  {32'hc5446c44, 32'h00000000} /* (23, 8, 0) {real, imag} */,
  {32'hc5485fc9, 32'h44db29a6} /* (23, 7, 31) {real, imag} */,
  {32'h446f3921, 32'hc3cb0544} /* (23, 7, 30) {real, imag} */,
  {32'h42c91dbe, 32'hc2bbfd38} /* (23, 7, 29) {real, imag} */,
  {32'hc2f16274, 32'hc1d75dce} /* (23, 7, 28) {real, imag} */,
  {32'h4309a334, 32'hc2e46984} /* (23, 7, 27) {real, imag} */,
  {32'h42702da6, 32'hc2cc1636} /* (23, 7, 26) {real, imag} */,
  {32'hc2cb581e, 32'h41db7b2d} /* (23, 7, 25) {real, imag} */,
  {32'h42edb8ec, 32'h418f2c16} /* (23, 7, 24) {real, imag} */,
  {32'h42b17c80, 32'hbfd53080} /* (23, 7, 23) {real, imag} */,
  {32'h4124d5e1, 32'h428b2079} /* (23, 7, 22) {real, imag} */,
  {32'hc22d6217, 32'h4035a340} /* (23, 7, 21) {real, imag} */,
  {32'h42ad6600, 32'h418f8e1a} /* (23, 7, 20) {real, imag} */,
  {32'h413f0f7c, 32'hc2815748} /* (23, 7, 19) {real, imag} */,
  {32'h421c745f, 32'h41aca27e} /* (23, 7, 18) {real, imag} */,
  {32'h4089d364, 32'h429b9c26} /* (23, 7, 17) {real, imag} */,
  {32'hc22adc6c, 32'h00000000} /* (23, 7, 16) {real, imag} */,
  {32'h4089d364, 32'hc29b9c26} /* (23, 7, 15) {real, imag} */,
  {32'h421c745f, 32'hc1aca27e} /* (23, 7, 14) {real, imag} */,
  {32'h413f0f7c, 32'h42815748} /* (23, 7, 13) {real, imag} */,
  {32'h42ad6600, 32'hc18f8e1a} /* (23, 7, 12) {real, imag} */,
  {32'hc22d6217, 32'hc035a340} /* (23, 7, 11) {real, imag} */,
  {32'h4124d5e1, 32'hc28b2079} /* (23, 7, 10) {real, imag} */,
  {32'h42b17c80, 32'h3fd53080} /* (23, 7, 9) {real, imag} */,
  {32'h42edb8ec, 32'hc18f2c16} /* (23, 7, 8) {real, imag} */,
  {32'hc2cb581e, 32'hc1db7b2d} /* (23, 7, 7) {real, imag} */,
  {32'h42702da6, 32'h42cc1636} /* (23, 7, 6) {real, imag} */,
  {32'h4309a334, 32'h42e46984} /* (23, 7, 5) {real, imag} */,
  {32'hc2f16274, 32'h41d75dce} /* (23, 7, 4) {real, imag} */,
  {32'h42c91dbe, 32'h42bbfd38} /* (23, 7, 3) {real, imag} */,
  {32'h446f3921, 32'h43cb0544} /* (23, 7, 2) {real, imag} */,
  {32'hc5485fc9, 32'hc4db29a6} /* (23, 7, 1) {real, imag} */,
  {32'hc56df3f4, 32'h00000000} /* (23, 7, 0) {real, imag} */,
  {32'hc5543844, 32'h450b3ef6} /* (23, 6, 31) {real, imag} */,
  {32'h443ea0fb, 32'hc417c97a} /* (23, 6, 30) {real, imag} */,
  {32'h4238c9a2, 32'h425cbc2d} /* (23, 6, 29) {real, imag} */,
  {32'hc2fc44c2, 32'h41df9b3a} /* (23, 6, 28) {real, imag} */,
  {32'h42fa863e, 32'hc2d403cb} /* (23, 6, 27) {real, imag} */,
  {32'hc136d3a3, 32'hc169003e} /* (23, 6, 26) {real, imag} */,
  {32'hc2979839, 32'hc17ad7b8} /* (23, 6, 25) {real, imag} */,
  {32'h42631a81, 32'hc275a252} /* (23, 6, 24) {real, imag} */,
  {32'hc0d4d838, 32'h40b27d24} /* (23, 6, 23) {real, imag} */,
  {32'hc27f8c48, 32'h420d22a0} /* (23, 6, 22) {real, imag} */,
  {32'hc2264d45, 32'hc2684e89} /* (23, 6, 21) {real, imag} */,
  {32'h41878788, 32'hc0b21ba0} /* (23, 6, 20) {real, imag} */,
  {32'hc214f676, 32'hc0dbc55c} /* (23, 6, 19) {real, imag} */,
  {32'h420a10ac, 32'hc1024066} /* (23, 6, 18) {real, imag} */,
  {32'hc1c702fb, 32'h41f44754} /* (23, 6, 17) {real, imag} */,
  {32'hc1f430c7, 32'h00000000} /* (23, 6, 16) {real, imag} */,
  {32'hc1c702fb, 32'hc1f44754} /* (23, 6, 15) {real, imag} */,
  {32'h420a10ac, 32'h41024066} /* (23, 6, 14) {real, imag} */,
  {32'hc214f676, 32'h40dbc55c} /* (23, 6, 13) {real, imag} */,
  {32'h41878788, 32'h40b21ba0} /* (23, 6, 12) {real, imag} */,
  {32'hc2264d45, 32'h42684e89} /* (23, 6, 11) {real, imag} */,
  {32'hc27f8c48, 32'hc20d22a0} /* (23, 6, 10) {real, imag} */,
  {32'hc0d4d838, 32'hc0b27d24} /* (23, 6, 9) {real, imag} */,
  {32'h42631a81, 32'h4275a252} /* (23, 6, 8) {real, imag} */,
  {32'hc2979839, 32'h417ad7b8} /* (23, 6, 7) {real, imag} */,
  {32'hc136d3a3, 32'h4169003e} /* (23, 6, 6) {real, imag} */,
  {32'h42fa863e, 32'h42d403cb} /* (23, 6, 5) {real, imag} */,
  {32'hc2fc44c2, 32'hc1df9b3a} /* (23, 6, 4) {real, imag} */,
  {32'h4238c9a2, 32'hc25cbc2d} /* (23, 6, 3) {real, imag} */,
  {32'h443ea0fb, 32'h4417c97a} /* (23, 6, 2) {real, imag} */,
  {32'hc5543844, 32'hc50b3ef6} /* (23, 6, 1) {real, imag} */,
  {32'hc5810825, 32'h00000000} /* (23, 6, 0) {real, imag} */,
  {32'hc54c8eeb, 32'h4538d601} /* (23, 5, 31) {real, imag} */,
  {32'h43675b68, 32'hc42c2312} /* (23, 5, 30) {real, imag} */,
  {32'h42d822fa, 32'hc1bc0a9c} /* (23, 5, 29) {real, imag} */,
  {32'h41b17936, 32'hc268171f} /* (23, 5, 28) {real, imag} */,
  {32'h4308380c, 32'h41ab0a38} /* (23, 5, 27) {real, imag} */,
  {32'hc16f22c2, 32'hc1e6a824} /* (23, 5, 26) {real, imag} */,
  {32'h4187a3a0, 32'h3f312500} /* (23, 5, 25) {real, imag} */,
  {32'hc28ff56a, 32'h41261c8d} /* (23, 5, 24) {real, imag} */,
  {32'h41c56b88, 32'hc2075910} /* (23, 5, 23) {real, imag} */,
  {32'hc2bf54e2, 32'hc208eafa} /* (23, 5, 22) {real, imag} */,
  {32'h421af306, 32'hc1eea3c9} /* (23, 5, 21) {real, imag} */,
  {32'h402be9ec, 32'h429894ee} /* (23, 5, 20) {real, imag} */,
  {32'hc1c303b4, 32'h420dd1ab} /* (23, 5, 19) {real, imag} */,
  {32'h41033a78, 32'hc20aea1c} /* (23, 5, 18) {real, imag} */,
  {32'h4262489e, 32'hc2502641} /* (23, 5, 17) {real, imag} */,
  {32'h40840208, 32'h00000000} /* (23, 5, 16) {real, imag} */,
  {32'h4262489e, 32'h42502641} /* (23, 5, 15) {real, imag} */,
  {32'h41033a78, 32'h420aea1c} /* (23, 5, 14) {real, imag} */,
  {32'hc1c303b4, 32'hc20dd1ab} /* (23, 5, 13) {real, imag} */,
  {32'h402be9ec, 32'hc29894ee} /* (23, 5, 12) {real, imag} */,
  {32'h421af306, 32'h41eea3c9} /* (23, 5, 11) {real, imag} */,
  {32'hc2bf54e2, 32'h4208eafa} /* (23, 5, 10) {real, imag} */,
  {32'h41c56b88, 32'h42075910} /* (23, 5, 9) {real, imag} */,
  {32'hc28ff56a, 32'hc1261c8d} /* (23, 5, 8) {real, imag} */,
  {32'h4187a3a0, 32'hbf312500} /* (23, 5, 7) {real, imag} */,
  {32'hc16f22c2, 32'h41e6a824} /* (23, 5, 6) {real, imag} */,
  {32'h4308380c, 32'hc1ab0a38} /* (23, 5, 5) {real, imag} */,
  {32'h41b17936, 32'h4268171f} /* (23, 5, 4) {real, imag} */,
  {32'h42d822fa, 32'h41bc0a9c} /* (23, 5, 3) {real, imag} */,
  {32'h43675b68, 32'h442c2312} /* (23, 5, 2) {real, imag} */,
  {32'hc54c8eeb, 32'hc538d601} /* (23, 5, 1) {real, imag} */,
  {32'hc5914ed7, 32'h00000000} /* (23, 5, 0) {real, imag} */,
  {32'hc5463803, 32'h455c3d95} /* (23, 4, 31) {real, imag} */,
  {32'hc28c95f0, 32'hc42ffb0e} /* (23, 4, 30) {real, imag} */,
  {32'h43116c9c, 32'hc302d2ef} /* (23, 4, 29) {real, imag} */,
  {32'h4308d1ef, 32'hc35328a2} /* (23, 4, 28) {real, imag} */,
  {32'h433fb7a6, 32'h4319233e} /* (23, 4, 27) {real, imag} */,
  {32'h42e380a6, 32'h4303b274} /* (23, 4, 26) {real, imag} */,
  {32'h42c2e41e, 32'hbf465280} /* (23, 4, 25) {real, imag} */,
  {32'hc2b2ffbf, 32'h418484b0} /* (23, 4, 24) {real, imag} */,
  {32'h42213677, 32'hc2856a3e} /* (23, 4, 23) {real, imag} */,
  {32'h422c2ee0, 32'hc276975a} /* (23, 4, 22) {real, imag} */,
  {32'h41c64808, 32'h4285cd83} /* (23, 4, 21) {real, imag} */,
  {32'h40c01d66, 32'hc2dc4ff0} /* (23, 4, 20) {real, imag} */,
  {32'hc20cb715, 32'h41ad930a} /* (23, 4, 19) {real, imag} */,
  {32'h406d05a0, 32'hc21f2f5c} /* (23, 4, 18) {real, imag} */,
  {32'h41d7f242, 32'hc2599b9c} /* (23, 4, 17) {real, imag} */,
  {32'hc147e9f8, 32'h00000000} /* (23, 4, 16) {real, imag} */,
  {32'h41d7f242, 32'h42599b9c} /* (23, 4, 15) {real, imag} */,
  {32'h406d05a0, 32'h421f2f5c} /* (23, 4, 14) {real, imag} */,
  {32'hc20cb715, 32'hc1ad930a} /* (23, 4, 13) {real, imag} */,
  {32'h40c01d66, 32'h42dc4ff0} /* (23, 4, 12) {real, imag} */,
  {32'h41c64808, 32'hc285cd83} /* (23, 4, 11) {real, imag} */,
  {32'h422c2ee0, 32'h4276975a} /* (23, 4, 10) {real, imag} */,
  {32'h42213677, 32'h42856a3e} /* (23, 4, 9) {real, imag} */,
  {32'hc2b2ffbf, 32'hc18484b0} /* (23, 4, 8) {real, imag} */,
  {32'h42c2e41e, 32'h3f465280} /* (23, 4, 7) {real, imag} */,
  {32'h42e380a6, 32'hc303b274} /* (23, 4, 6) {real, imag} */,
  {32'h433fb7a6, 32'hc319233e} /* (23, 4, 5) {real, imag} */,
  {32'h4308d1ef, 32'h435328a2} /* (23, 4, 4) {real, imag} */,
  {32'h43116c9c, 32'h4302d2ef} /* (23, 4, 3) {real, imag} */,
  {32'hc28c95f0, 32'h442ffb0e} /* (23, 4, 2) {real, imag} */,
  {32'hc5463803, 32'hc55c3d95} /* (23, 4, 1) {real, imag} */,
  {32'hc59cc802, 32'h00000000} /* (23, 4, 0) {real, imag} */,
  {32'hc54b27fd, 32'h45631154} /* (23, 3, 31) {real, imag} */,
  {32'hc3bab94a, 32'hc45c0adf} /* (23, 3, 30) {real, imag} */,
  {32'h42f70486, 32'h4106a898} /* (23, 3, 29) {real, imag} */,
  {32'h426929fe, 32'hc39df64f} /* (23, 3, 28) {real, imag} */,
  {32'h436b9ec5, 32'h43135c7d} /* (23, 3, 27) {real, imag} */,
  {32'h430a179a, 32'h4173140c} /* (23, 3, 26) {real, imag} */,
  {32'h42337533, 32'h4305bd04} /* (23, 3, 25) {real, imag} */,
  {32'hc2434851, 32'hc22c80d8} /* (23, 3, 24) {real, imag} */,
  {32'h4295c05a, 32'hc1c90673} /* (23, 3, 23) {real, imag} */,
  {32'h40d39e28, 32'h409d1660} /* (23, 3, 22) {real, imag} */,
  {32'h4223639a, 32'hc1fd7728} /* (23, 3, 21) {real, imag} */,
  {32'hc1d14d57, 32'h3fb72168} /* (23, 3, 20) {real, imag} */,
  {32'h413a7390, 32'hc284ffd2} /* (23, 3, 19) {real, imag} */,
  {32'hc2de51b6, 32'h428ef7d4} /* (23, 3, 18) {real, imag} */,
  {32'hc1ef2eb1, 32'hc1f5f0d5} /* (23, 3, 17) {real, imag} */,
  {32'hc31f5d9a, 32'h00000000} /* (23, 3, 16) {real, imag} */,
  {32'hc1ef2eb1, 32'h41f5f0d5} /* (23, 3, 15) {real, imag} */,
  {32'hc2de51b6, 32'hc28ef7d4} /* (23, 3, 14) {real, imag} */,
  {32'h413a7390, 32'h4284ffd2} /* (23, 3, 13) {real, imag} */,
  {32'hc1d14d57, 32'hbfb72168} /* (23, 3, 12) {real, imag} */,
  {32'h4223639a, 32'h41fd7728} /* (23, 3, 11) {real, imag} */,
  {32'h40d39e28, 32'hc09d1660} /* (23, 3, 10) {real, imag} */,
  {32'h4295c05a, 32'h41c90673} /* (23, 3, 9) {real, imag} */,
  {32'hc2434851, 32'h422c80d8} /* (23, 3, 8) {real, imag} */,
  {32'h42337533, 32'hc305bd04} /* (23, 3, 7) {real, imag} */,
  {32'h430a179a, 32'hc173140c} /* (23, 3, 6) {real, imag} */,
  {32'h436b9ec5, 32'hc3135c7d} /* (23, 3, 5) {real, imag} */,
  {32'h426929fe, 32'h439df64f} /* (23, 3, 4) {real, imag} */,
  {32'h42f70486, 32'hc106a898} /* (23, 3, 3) {real, imag} */,
  {32'hc3bab94a, 32'h445c0adf} /* (23, 3, 2) {real, imag} */,
  {32'hc54b27fd, 32'hc5631154} /* (23, 3, 1) {real, imag} */,
  {32'hc59e39b4, 32'h00000000} /* (23, 3, 0) {real, imag} */,
  {32'hc53f4755, 32'h456401f6} /* (23, 2, 31) {real, imag} */,
  {32'hc384ec55, 32'hc4564150} /* (23, 2, 30) {real, imag} */,
  {32'h435e3f74, 32'h4101f212} /* (23, 2, 29) {real, imag} */,
  {32'h42238cf8, 32'hc3b2d2a4} /* (23, 2, 28) {real, imag} */,
  {32'h439a624b, 32'hc1cfb150} /* (23, 2, 27) {real, imag} */,
  {32'hc2002c8c, 32'h410e8060} /* (23, 2, 26) {real, imag} */,
  {32'h428f230e, 32'h42ce2692} /* (23, 2, 25) {real, imag} */,
  {32'hc2d26c96, 32'h40e14d58} /* (23, 2, 24) {real, imag} */,
  {32'hc170cb9e, 32'hc2e83dfa} /* (23, 2, 23) {real, imag} */,
  {32'hc2892f04, 32'h42aefe5e} /* (23, 2, 22) {real, imag} */,
  {32'h42a488d3, 32'h4242097c} /* (23, 2, 21) {real, imag} */,
  {32'h3f5ffe80, 32'h43022782} /* (23, 2, 20) {real, imag} */,
  {32'hc29812b4, 32'h42cec2d0} /* (23, 2, 19) {real, imag} */,
  {32'h3fcfa1a0, 32'hc262768a} /* (23, 2, 18) {real, imag} */,
  {32'h420f46e7, 32'hc25f5ade} /* (23, 2, 17) {real, imag} */,
  {32'hc28452b6, 32'h00000000} /* (23, 2, 16) {real, imag} */,
  {32'h420f46e7, 32'h425f5ade} /* (23, 2, 15) {real, imag} */,
  {32'h3fcfa1a0, 32'h4262768a} /* (23, 2, 14) {real, imag} */,
  {32'hc29812b4, 32'hc2cec2d0} /* (23, 2, 13) {real, imag} */,
  {32'h3f5ffe80, 32'hc3022782} /* (23, 2, 12) {real, imag} */,
  {32'h42a488d3, 32'hc242097c} /* (23, 2, 11) {real, imag} */,
  {32'hc2892f04, 32'hc2aefe5e} /* (23, 2, 10) {real, imag} */,
  {32'hc170cb9e, 32'h42e83dfa} /* (23, 2, 9) {real, imag} */,
  {32'hc2d26c96, 32'hc0e14d58} /* (23, 2, 8) {real, imag} */,
  {32'h428f230e, 32'hc2ce2692} /* (23, 2, 7) {real, imag} */,
  {32'hc2002c8c, 32'hc10e8060} /* (23, 2, 6) {real, imag} */,
  {32'h439a624b, 32'h41cfb150} /* (23, 2, 5) {real, imag} */,
  {32'h42238cf8, 32'h43b2d2a4} /* (23, 2, 4) {real, imag} */,
  {32'h435e3f74, 32'hc101f212} /* (23, 2, 3) {real, imag} */,
  {32'hc384ec55, 32'h44564150} /* (23, 2, 2) {real, imag} */,
  {32'hc53f4755, 32'hc56401f6} /* (23, 2, 1) {real, imag} */,
  {32'hc5a4b13c, 32'h00000000} /* (23, 2, 0) {real, imag} */,
  {32'hc543445e, 32'h45537ada} /* (23, 1, 31) {real, imag} */,
  {32'hc317e736, 32'hc425f07e} /* (23, 1, 30) {real, imag} */,
  {32'h439e758e, 32'hc210d2b2} /* (23, 1, 29) {real, imag} */,
  {32'h42ae3520, 32'hc39d918e} /* (23, 1, 28) {real, imag} */,
  {32'h435f1122, 32'h4266febe} /* (23, 1, 27) {real, imag} */,
  {32'hc2d617c7, 32'h42377366} /* (23, 1, 26) {real, imag} */,
  {32'hc1f281fc, 32'hc114f8d0} /* (23, 1, 25) {real, imag} */,
  {32'h41c7c2d0, 32'hc058eff8} /* (23, 1, 24) {real, imag} */,
  {32'h4243d84e, 32'h4203f198} /* (23, 1, 23) {real, imag} */,
  {32'hc2a02d57, 32'hc2d87cca} /* (23, 1, 22) {real, imag} */,
  {32'h4274bfdc, 32'hc234210c} /* (23, 1, 21) {real, imag} */,
  {32'hc23f925a, 32'h421231ec} /* (23, 1, 20) {real, imag} */,
  {32'hc2498c42, 32'h41f2cb02} /* (23, 1, 19) {real, imag} */,
  {32'hc1bf0533, 32'hc1c4c636} /* (23, 1, 18) {real, imag} */,
  {32'h42968a65, 32'hc247b14c} /* (23, 1, 17) {real, imag} */,
  {32'h42925085, 32'h00000000} /* (23, 1, 16) {real, imag} */,
  {32'h42968a65, 32'h4247b14c} /* (23, 1, 15) {real, imag} */,
  {32'hc1bf0533, 32'h41c4c636} /* (23, 1, 14) {real, imag} */,
  {32'hc2498c42, 32'hc1f2cb02} /* (23, 1, 13) {real, imag} */,
  {32'hc23f925a, 32'hc21231ec} /* (23, 1, 12) {real, imag} */,
  {32'h4274bfdc, 32'h4234210c} /* (23, 1, 11) {real, imag} */,
  {32'hc2a02d57, 32'h42d87cca} /* (23, 1, 10) {real, imag} */,
  {32'h4243d84e, 32'hc203f198} /* (23, 1, 9) {real, imag} */,
  {32'h41c7c2d0, 32'h4058eff8} /* (23, 1, 8) {real, imag} */,
  {32'hc1f281fc, 32'h4114f8d0} /* (23, 1, 7) {real, imag} */,
  {32'hc2d617c7, 32'hc2377366} /* (23, 1, 6) {real, imag} */,
  {32'h435f1122, 32'hc266febe} /* (23, 1, 5) {real, imag} */,
  {32'h42ae3520, 32'h439d918e} /* (23, 1, 4) {real, imag} */,
  {32'h439e758e, 32'h4210d2b2} /* (23, 1, 3) {real, imag} */,
  {32'hc317e736, 32'h4425f07e} /* (23, 1, 2) {real, imag} */,
  {32'hc543445e, 32'hc5537ada} /* (23, 1, 1) {real, imag} */,
  {32'hc59860d5, 32'h00000000} /* (23, 1, 0) {real, imag} */,
  {32'hc54ce74e, 32'h452c21bf} /* (23, 0, 31) {real, imag} */,
  {32'h43565a38, 32'hc3e30377} /* (23, 0, 30) {real, imag} */,
  {32'h430ea3bf, 32'hc13d9fd4} /* (23, 0, 29) {real, imag} */,
  {32'h428bb0c8, 32'hc365a2cc} /* (23, 0, 28) {real, imag} */,
  {32'h4233790c, 32'h42b7502b} /* (23, 0, 27) {real, imag} */,
  {32'hbfdbf280, 32'hc2185360} /* (23, 0, 26) {real, imag} */,
  {32'h42003b10, 32'h40a1d0b8} /* (23, 0, 25) {real, imag} */,
  {32'h4205e2ed, 32'h41998b76} /* (23, 0, 24) {real, imag} */,
  {32'h4292c37c, 32'h42683f9a} /* (23, 0, 23) {real, imag} */,
  {32'h3ebcf6b0, 32'hc2be6e5a} /* (23, 0, 22) {real, imag} */,
  {32'hc29cffce, 32'hc21eff03} /* (23, 0, 21) {real, imag} */,
  {32'h41b94a76, 32'h418832dc} /* (23, 0, 20) {real, imag} */,
  {32'h40887912, 32'h420ca853} /* (23, 0, 19) {real, imag} */,
  {32'hc23188ea, 32'h4207139c} /* (23, 0, 18) {real, imag} */,
  {32'h4189195d, 32'hc260fc60} /* (23, 0, 17) {real, imag} */,
  {32'h426814a8, 32'h00000000} /* (23, 0, 16) {real, imag} */,
  {32'h4189195d, 32'h4260fc60} /* (23, 0, 15) {real, imag} */,
  {32'hc23188ea, 32'hc207139c} /* (23, 0, 14) {real, imag} */,
  {32'h40887912, 32'hc20ca853} /* (23, 0, 13) {real, imag} */,
  {32'h41b94a76, 32'hc18832dc} /* (23, 0, 12) {real, imag} */,
  {32'hc29cffce, 32'h421eff03} /* (23, 0, 11) {real, imag} */,
  {32'h3ebcf6b0, 32'h42be6e5a} /* (23, 0, 10) {real, imag} */,
  {32'h4292c37c, 32'hc2683f9a} /* (23, 0, 9) {real, imag} */,
  {32'h4205e2ed, 32'hc1998b76} /* (23, 0, 8) {real, imag} */,
  {32'h42003b10, 32'hc0a1d0b8} /* (23, 0, 7) {real, imag} */,
  {32'hbfdbf280, 32'h42185360} /* (23, 0, 6) {real, imag} */,
  {32'h4233790c, 32'hc2b7502b} /* (23, 0, 5) {real, imag} */,
  {32'h428bb0c8, 32'h4365a2cc} /* (23, 0, 4) {real, imag} */,
  {32'h430ea3bf, 32'h413d9fd4} /* (23, 0, 3) {real, imag} */,
  {32'h43565a38, 32'h43e30377} /* (23, 0, 2) {real, imag} */,
  {32'hc54ce74e, 32'hc52c21bf} /* (23, 0, 1) {real, imag} */,
  {32'hc5967900, 32'h00000000} /* (23, 0, 0) {real, imag} */,
  {32'hc57d526d, 32'h45153968} /* (22, 31, 31) {real, imag} */,
  {32'h443c123b, 32'hc3dce955} /* (22, 31, 30) {real, imag} */,
  {32'h41b07878, 32'h41bf9e88} /* (22, 31, 29) {real, imag} */,
  {32'hc2efaa3a, 32'hc1e035f8} /* (22, 31, 28) {real, imag} */,
  {32'h42be0aa6, 32'hc1bc9630} /* (22, 31, 27) {real, imag} */,
  {32'h42205888, 32'hc1735a26} /* (22, 31, 26) {real, imag} */,
  {32'hc24fca44, 32'h41b65660} /* (22, 31, 25) {real, imag} */,
  {32'hc0a72e34, 32'hc2592186} /* (22, 31, 24) {real, imag} */,
  {32'h3febc888, 32'h41d8b79a} /* (22, 31, 23) {real, imag} */,
  {32'h42c8b8ac, 32'hc256b8bc} /* (22, 31, 22) {real, imag} */,
  {32'h4203bc4c, 32'hbf5302e0} /* (22, 31, 21) {real, imag} */,
  {32'hc1fbf2a1, 32'hc28a1b70} /* (22, 31, 20) {real, imag} */,
  {32'h42568739, 32'h424e8e96} /* (22, 31, 19) {real, imag} */,
  {32'h4205ee50, 32'h4138cb36} /* (22, 31, 18) {real, imag} */,
  {32'hc10e1496, 32'h40b63462} /* (22, 31, 17) {real, imag} */,
  {32'h40d557e6, 32'h00000000} /* (22, 31, 16) {real, imag} */,
  {32'hc10e1496, 32'hc0b63462} /* (22, 31, 15) {real, imag} */,
  {32'h4205ee50, 32'hc138cb36} /* (22, 31, 14) {real, imag} */,
  {32'h42568739, 32'hc24e8e96} /* (22, 31, 13) {real, imag} */,
  {32'hc1fbf2a1, 32'h428a1b70} /* (22, 31, 12) {real, imag} */,
  {32'h4203bc4c, 32'h3f5302e0} /* (22, 31, 11) {real, imag} */,
  {32'h42c8b8ac, 32'h4256b8bc} /* (22, 31, 10) {real, imag} */,
  {32'h3febc888, 32'hc1d8b79a} /* (22, 31, 9) {real, imag} */,
  {32'hc0a72e34, 32'h42592186} /* (22, 31, 8) {real, imag} */,
  {32'hc24fca44, 32'hc1b65660} /* (22, 31, 7) {real, imag} */,
  {32'h42205888, 32'h41735a26} /* (22, 31, 6) {real, imag} */,
  {32'h42be0aa6, 32'h41bc9630} /* (22, 31, 5) {real, imag} */,
  {32'hc2efaa3a, 32'h41e035f8} /* (22, 31, 4) {real, imag} */,
  {32'h41b07878, 32'hc1bf9e88} /* (22, 31, 3) {real, imag} */,
  {32'h443c123b, 32'h43dce955} /* (22, 31, 2) {real, imag} */,
  {32'hc57d526d, 32'hc5153968} /* (22, 31, 1) {real, imag} */,
  {32'hc5a381fb, 32'h00000000} /* (22, 31, 0) {real, imag} */,
  {32'hc58fe08b, 32'h44fb98f6} /* (22, 30, 31) {real, imag} */,
  {32'h449c5391, 32'hc3c3e39c} /* (22, 30, 30) {real, imag} */,
  {32'hc20599ea, 32'hc1b83612} /* (22, 30, 29) {real, imag} */,
  {32'hc39fce2d, 32'h41881eb0} /* (22, 30, 28) {real, imag} */,
  {32'h436c2e92, 32'h420d6cbe} /* (22, 30, 27) {real, imag} */,
  {32'h421293e1, 32'hc0a23d40} /* (22, 30, 26) {real, imag} */,
  {32'hc2744db7, 32'hc28f8763} /* (22, 30, 25) {real, imag} */,
  {32'h41f119d0, 32'hc2b0686f} /* (22, 30, 24) {real, imag} */,
  {32'hc3024fcf, 32'hc20b003c} /* (22, 30, 23) {real, imag} */,
  {32'h42a5f1e2, 32'h41da5a7e} /* (22, 30, 22) {real, imag} */,
  {32'h42a5e53f, 32'h41a901f8} /* (22, 30, 21) {real, imag} */,
  {32'hc28be628, 32'h419a224e} /* (22, 30, 20) {real, imag} */,
  {32'h4213ce5c, 32'h4277e912} /* (22, 30, 19) {real, imag} */,
  {32'h41e7bb7f, 32'hc2c9b0da} /* (22, 30, 18) {real, imag} */,
  {32'hc1fd60c9, 32'hc1f7593e} /* (22, 30, 17) {real, imag} */,
  {32'h424eac42, 32'h00000000} /* (22, 30, 16) {real, imag} */,
  {32'hc1fd60c9, 32'h41f7593e} /* (22, 30, 15) {real, imag} */,
  {32'h41e7bb7f, 32'h42c9b0da} /* (22, 30, 14) {real, imag} */,
  {32'h4213ce5c, 32'hc277e912} /* (22, 30, 13) {real, imag} */,
  {32'hc28be628, 32'hc19a224e} /* (22, 30, 12) {real, imag} */,
  {32'h42a5e53f, 32'hc1a901f8} /* (22, 30, 11) {real, imag} */,
  {32'h42a5f1e2, 32'hc1da5a7e} /* (22, 30, 10) {real, imag} */,
  {32'hc3024fcf, 32'h420b003c} /* (22, 30, 9) {real, imag} */,
  {32'h41f119d0, 32'h42b0686f} /* (22, 30, 8) {real, imag} */,
  {32'hc2744db7, 32'h428f8763} /* (22, 30, 7) {real, imag} */,
  {32'h421293e1, 32'h40a23d40} /* (22, 30, 6) {real, imag} */,
  {32'h436c2e92, 32'hc20d6cbe} /* (22, 30, 5) {real, imag} */,
  {32'hc39fce2d, 32'hc1881eb0} /* (22, 30, 4) {real, imag} */,
  {32'hc20599ea, 32'h41b83612} /* (22, 30, 3) {real, imag} */,
  {32'h449c5391, 32'h43c3e39c} /* (22, 30, 2) {real, imag} */,
  {32'hc58fe08b, 32'hc4fb98f6} /* (22, 30, 1) {real, imag} */,
  {32'hc5ab546d, 32'h00000000} /* (22, 30, 0) {real, imag} */,
  {32'hc59db42a, 32'h44cba777} /* (22, 29, 31) {real, imag} */,
  {32'h44c401aa, 32'hc3b2acc2} /* (22, 29, 30) {real, imag} */,
  {32'hc2b68426, 32'hc2616c00} /* (22, 29, 29) {real, imag} */,
  {32'hc385da77, 32'h42c63643} /* (22, 29, 28) {real, imag} */,
  {32'h434ae450, 32'hc35e9cdf} /* (22, 29, 27) {real, imag} */,
  {32'hc2809994, 32'hc2659a61} /* (22, 29, 26) {real, imag} */,
  {32'hc260b0bb, 32'hc227730a} /* (22, 29, 25) {real, imag} */,
  {32'h426d6d5c, 32'hc33012c8} /* (22, 29, 24) {real, imag} */,
  {32'hc22284e2, 32'hc13d5c16} /* (22, 29, 23) {real, imag} */,
  {32'h430b15ac, 32'hc1db9f74} /* (22, 29, 22) {real, imag} */,
  {32'h41ebd520, 32'hc251f742} /* (22, 29, 21) {real, imag} */,
  {32'h418248f0, 32'h42668e88} /* (22, 29, 20) {real, imag} */,
  {32'h41811a5a, 32'hc2c83984} /* (22, 29, 19) {real, imag} */,
  {32'hc1c9f636, 32'h423b3de2} /* (22, 29, 18) {real, imag} */,
  {32'h41bdefe4, 32'h41f329a7} /* (22, 29, 17) {real, imag} */,
  {32'hc0f48888, 32'h00000000} /* (22, 29, 16) {real, imag} */,
  {32'h41bdefe4, 32'hc1f329a7} /* (22, 29, 15) {real, imag} */,
  {32'hc1c9f636, 32'hc23b3de2} /* (22, 29, 14) {real, imag} */,
  {32'h41811a5a, 32'h42c83984} /* (22, 29, 13) {real, imag} */,
  {32'h418248f0, 32'hc2668e88} /* (22, 29, 12) {real, imag} */,
  {32'h41ebd520, 32'h4251f742} /* (22, 29, 11) {real, imag} */,
  {32'h430b15ac, 32'h41db9f74} /* (22, 29, 10) {real, imag} */,
  {32'hc22284e2, 32'h413d5c16} /* (22, 29, 9) {real, imag} */,
  {32'h426d6d5c, 32'h433012c8} /* (22, 29, 8) {real, imag} */,
  {32'hc260b0bb, 32'h4227730a} /* (22, 29, 7) {real, imag} */,
  {32'hc2809994, 32'h42659a61} /* (22, 29, 6) {real, imag} */,
  {32'h434ae450, 32'h435e9cdf} /* (22, 29, 5) {real, imag} */,
  {32'hc385da77, 32'hc2c63643} /* (22, 29, 4) {real, imag} */,
  {32'hc2b68426, 32'h42616c00} /* (22, 29, 3) {real, imag} */,
  {32'h44c401aa, 32'h43b2acc2} /* (22, 29, 2) {real, imag} */,
  {32'hc59db42a, 32'hc4cba777} /* (22, 29, 1) {real, imag} */,
  {32'hc5abf71c, 32'h00000000} /* (22, 29, 0) {real, imag} */,
  {32'hc5a58dc3, 32'h44aa7dc2} /* (22, 28, 31) {real, imag} */,
  {32'h44e691e8, 32'hc3b34409} /* (22, 28, 30) {real, imag} */,
  {32'hc21b0fcc, 32'hc2e55dd0} /* (22, 28, 29) {real, imag} */,
  {32'hc35d97aa, 32'h432d0bef} /* (22, 28, 28) {real, imag} */,
  {32'h437467eb, 32'hc305d509} /* (22, 28, 27) {real, imag} */,
  {32'hc04e51f0, 32'hc28a947b} /* (22, 28, 26) {real, imag} */,
  {32'hc0b85e8c, 32'h4287858c} /* (22, 28, 25) {real, imag} */,
  {32'h427fc589, 32'hc349ca06} /* (22, 28, 24) {real, imag} */,
  {32'h411b8ea4, 32'h428ce0b4} /* (22, 28, 23) {real, imag} */,
  {32'h41023cde, 32'hc0dff778} /* (22, 28, 22) {real, imag} */,
  {32'h424ee2f4, 32'h428df3cb} /* (22, 28, 21) {real, imag} */,
  {32'hc1b81076, 32'hc26d24df} /* (22, 28, 20) {real, imag} */,
  {32'hc1fcd356, 32'h41fa4876} /* (22, 28, 19) {real, imag} */,
  {32'h418161b6, 32'h421534ad} /* (22, 28, 18) {real, imag} */,
  {32'h41a0e8ec, 32'h41bb54ba} /* (22, 28, 17) {real, imag} */,
  {32'h40fe0fcc, 32'h00000000} /* (22, 28, 16) {real, imag} */,
  {32'h41a0e8ec, 32'hc1bb54ba} /* (22, 28, 15) {real, imag} */,
  {32'h418161b6, 32'hc21534ad} /* (22, 28, 14) {real, imag} */,
  {32'hc1fcd356, 32'hc1fa4876} /* (22, 28, 13) {real, imag} */,
  {32'hc1b81076, 32'h426d24df} /* (22, 28, 12) {real, imag} */,
  {32'h424ee2f4, 32'hc28df3cb} /* (22, 28, 11) {real, imag} */,
  {32'h41023cde, 32'h40dff778} /* (22, 28, 10) {real, imag} */,
  {32'h411b8ea4, 32'hc28ce0b4} /* (22, 28, 9) {real, imag} */,
  {32'h427fc589, 32'h4349ca06} /* (22, 28, 8) {real, imag} */,
  {32'hc0b85e8c, 32'hc287858c} /* (22, 28, 7) {real, imag} */,
  {32'hc04e51f0, 32'h428a947b} /* (22, 28, 6) {real, imag} */,
  {32'h437467eb, 32'h4305d509} /* (22, 28, 5) {real, imag} */,
  {32'hc35d97aa, 32'hc32d0bef} /* (22, 28, 4) {real, imag} */,
  {32'hc21b0fcc, 32'h42e55dd0} /* (22, 28, 3) {real, imag} */,
  {32'h44e691e8, 32'h43b34409} /* (22, 28, 2) {real, imag} */,
  {32'hc5a58dc3, 32'hc4aa7dc2} /* (22, 28, 1) {real, imag} */,
  {32'hc5b0a1ab, 32'h00000000} /* (22, 28, 0) {real, imag} */,
  {32'hc5a5aa94, 32'h44750a72} /* (22, 27, 31) {real, imag} */,
  {32'h44ebd140, 32'hc3c66bda} /* (22, 27, 30) {real, imag} */,
  {32'h42a4d861, 32'hc196337c} /* (22, 27, 29) {real, imag} */,
  {32'hc359d8e7, 32'hc0e70d20} /* (22, 27, 28) {real, imag} */,
  {32'h43344539, 32'hc3293df4} /* (22, 27, 27) {real, imag} */,
  {32'hc1888096, 32'h4294f6ad} /* (22, 27, 26) {real, imag} */,
  {32'hc31acee0, 32'h428b1f80} /* (22, 27, 25) {real, imag} */,
  {32'hc29374f8, 32'hc20625a0} /* (22, 27, 24) {real, imag} */,
  {32'h4158b290, 32'hc2905754} /* (22, 27, 23) {real, imag} */,
  {32'h42b1311d, 32'h419ed4c8} /* (22, 27, 22) {real, imag} */,
  {32'h423484a8, 32'hc26659d5} /* (22, 27, 21) {real, imag} */,
  {32'hc291bed8, 32'hc25d3d1c} /* (22, 27, 20) {real, imag} */,
  {32'hc1c52a36, 32'h410c01c8} /* (22, 27, 19) {real, imag} */,
  {32'hc24d5d1e, 32'hc24e7878} /* (22, 27, 18) {real, imag} */,
  {32'h41cb7e88, 32'hc173ca80} /* (22, 27, 17) {real, imag} */,
  {32'h41229631, 32'h00000000} /* (22, 27, 16) {real, imag} */,
  {32'h41cb7e88, 32'h4173ca80} /* (22, 27, 15) {real, imag} */,
  {32'hc24d5d1e, 32'h424e7878} /* (22, 27, 14) {real, imag} */,
  {32'hc1c52a36, 32'hc10c01c8} /* (22, 27, 13) {real, imag} */,
  {32'hc291bed8, 32'h425d3d1c} /* (22, 27, 12) {real, imag} */,
  {32'h423484a8, 32'h426659d5} /* (22, 27, 11) {real, imag} */,
  {32'h42b1311d, 32'hc19ed4c8} /* (22, 27, 10) {real, imag} */,
  {32'h4158b290, 32'h42905754} /* (22, 27, 9) {real, imag} */,
  {32'hc29374f8, 32'h420625a0} /* (22, 27, 8) {real, imag} */,
  {32'hc31acee0, 32'hc28b1f80} /* (22, 27, 7) {real, imag} */,
  {32'hc1888096, 32'hc294f6ad} /* (22, 27, 6) {real, imag} */,
  {32'h43344539, 32'h43293df4} /* (22, 27, 5) {real, imag} */,
  {32'hc359d8e7, 32'h40e70d20} /* (22, 27, 4) {real, imag} */,
  {32'h42a4d861, 32'h4196337c} /* (22, 27, 3) {real, imag} */,
  {32'h44ebd140, 32'h43c66bda} /* (22, 27, 2) {real, imag} */,
  {32'hc5a5aa94, 32'hc4750a72} /* (22, 27, 1) {real, imag} */,
  {32'hc5b04050, 32'h00000000} /* (22, 27, 0) {real, imag} */,
  {32'hc59c964c, 32'h446ad84a} /* (22, 26, 31) {real, imag} */,
  {32'h44e6f03a, 32'hc3cf5658} /* (22, 26, 30) {real, imag} */,
  {32'hc10fd04a, 32'hc25daf91} /* (22, 26, 29) {real, imag} */,
  {32'hc3854caa, 32'hc0ec56d8} /* (22, 26, 28) {real, imag} */,
  {32'h439a8b5a, 32'hc35f8dc6} /* (22, 26, 27) {real, imag} */,
  {32'h4187ff04, 32'h428efa38} /* (22, 26, 26) {real, imag} */,
  {32'hc2b10d41, 32'hc21f6664} /* (22, 26, 25) {real, imag} */,
  {32'h420ebdb0, 32'hc27a4188} /* (22, 26, 24) {real, imag} */,
  {32'h41aecaac, 32'hc1cfd6ce} /* (22, 26, 23) {real, imag} */,
  {32'hc2030906, 32'h42c317a6} /* (22, 26, 22) {real, imag} */,
  {32'hc20f3682, 32'hc2f1e53c} /* (22, 26, 21) {real, imag} */,
  {32'h42ac5350, 32'hc24ed240} /* (22, 26, 20) {real, imag} */,
  {32'h422b28d8, 32'h419d13b3} /* (22, 26, 19) {real, imag} */,
  {32'h41d8e926, 32'h41ee81e8} /* (22, 26, 18) {real, imag} */,
  {32'h418d9736, 32'hc2013faf} /* (22, 26, 17) {real, imag} */,
  {32'hc17e1372, 32'h00000000} /* (22, 26, 16) {real, imag} */,
  {32'h418d9736, 32'h42013faf} /* (22, 26, 15) {real, imag} */,
  {32'h41d8e926, 32'hc1ee81e8} /* (22, 26, 14) {real, imag} */,
  {32'h422b28d8, 32'hc19d13b3} /* (22, 26, 13) {real, imag} */,
  {32'h42ac5350, 32'h424ed240} /* (22, 26, 12) {real, imag} */,
  {32'hc20f3682, 32'h42f1e53c} /* (22, 26, 11) {real, imag} */,
  {32'hc2030906, 32'hc2c317a6} /* (22, 26, 10) {real, imag} */,
  {32'h41aecaac, 32'h41cfd6ce} /* (22, 26, 9) {real, imag} */,
  {32'h420ebdb0, 32'h427a4188} /* (22, 26, 8) {real, imag} */,
  {32'hc2b10d41, 32'h421f6664} /* (22, 26, 7) {real, imag} */,
  {32'h4187ff04, 32'hc28efa38} /* (22, 26, 6) {real, imag} */,
  {32'h439a8b5a, 32'h435f8dc6} /* (22, 26, 5) {real, imag} */,
  {32'hc3854caa, 32'h40ec56d8} /* (22, 26, 4) {real, imag} */,
  {32'hc10fd04a, 32'h425daf91} /* (22, 26, 3) {real, imag} */,
  {32'h44e6f03a, 32'h43cf5658} /* (22, 26, 2) {real, imag} */,
  {32'hc59c964c, 32'hc46ad84a} /* (22, 26, 1) {real, imag} */,
  {32'hc5a993f6, 32'h00000000} /* (22, 26, 0) {real, imag} */,
  {32'hc592013c, 32'h443af51f} /* (22, 25, 31) {real, imag} */,
  {32'h44e85ea2, 32'hc3a75e27} /* (22, 25, 30) {real, imag} */,
  {32'hc306334c, 32'hc28bc1ca} /* (22, 25, 29) {real, imag} */,
  {32'hc3530d8f, 32'h42c30b82} /* (22, 25, 28) {real, imag} */,
  {32'h43816ce0, 32'hc2d6e804} /* (22, 25, 27) {real, imag} */,
  {32'h41d61536, 32'hc168f132} /* (22, 25, 26) {real, imag} */,
  {32'hc2b3c6ed, 32'hc244f47e} /* (22, 25, 25) {real, imag} */,
  {32'h42a1ce93, 32'hc282a0b4} /* (22, 25, 24) {real, imag} */,
  {32'h429a5438, 32'hc1df65e8} /* (22, 25, 23) {real, imag} */,
  {32'hbfd32aa0, 32'hc15588d8} /* (22, 25, 22) {real, imag} */,
  {32'hc209fad8, 32'hc236e3fb} /* (22, 25, 21) {real, imag} */,
  {32'hc166313d, 32'h426a5cfd} /* (22, 25, 20) {real, imag} */,
  {32'h423e1aae, 32'h409dd1f8} /* (22, 25, 19) {real, imag} */,
  {32'h42eee210, 32'hc1a0cae3} /* (22, 25, 18) {real, imag} */,
  {32'hc11f08c6, 32'h419f0b70} /* (22, 25, 17) {real, imag} */,
  {32'hc1e40055, 32'h00000000} /* (22, 25, 16) {real, imag} */,
  {32'hc11f08c6, 32'hc19f0b70} /* (22, 25, 15) {real, imag} */,
  {32'h42eee210, 32'h41a0cae3} /* (22, 25, 14) {real, imag} */,
  {32'h423e1aae, 32'hc09dd1f8} /* (22, 25, 13) {real, imag} */,
  {32'hc166313d, 32'hc26a5cfd} /* (22, 25, 12) {real, imag} */,
  {32'hc209fad8, 32'h4236e3fb} /* (22, 25, 11) {real, imag} */,
  {32'hbfd32aa0, 32'h415588d8} /* (22, 25, 10) {real, imag} */,
  {32'h429a5438, 32'h41df65e8} /* (22, 25, 9) {real, imag} */,
  {32'h42a1ce93, 32'h4282a0b4} /* (22, 25, 8) {real, imag} */,
  {32'hc2b3c6ed, 32'h4244f47e} /* (22, 25, 7) {real, imag} */,
  {32'h41d61536, 32'h4168f132} /* (22, 25, 6) {real, imag} */,
  {32'h43816ce0, 32'h42d6e804} /* (22, 25, 5) {real, imag} */,
  {32'hc3530d8f, 32'hc2c30b82} /* (22, 25, 4) {real, imag} */,
  {32'hc306334c, 32'h428bc1ca} /* (22, 25, 3) {real, imag} */,
  {32'h44e85ea2, 32'h43a75e27} /* (22, 25, 2) {real, imag} */,
  {32'hc592013c, 32'hc43af51f} /* (22, 25, 1) {real, imag} */,
  {32'hc59bd282, 32'h00000000} /* (22, 25, 0) {real, imag} */,
  {32'hc5848d57, 32'h440c892a} /* (22, 24, 31) {real, imag} */,
  {32'h44dd1d48, 32'hc3428386} /* (22, 24, 30) {real, imag} */,
  {32'hc2f992da, 32'h428ca6b5} /* (22, 24, 29) {real, imag} */,
  {32'hc22e04c8, 32'h43264515} /* (22, 24, 28) {real, imag} */,
  {32'h43501d60, 32'hc300e333} /* (22, 24, 27) {real, imag} */,
  {32'h423f7984, 32'hc20c71c7} /* (22, 24, 26) {real, imag} */,
  {32'h423bc214, 32'h42bbdd4e} /* (22, 24, 25) {real, imag} */,
  {32'h428bacf6, 32'hc23ae646} /* (22, 24, 24) {real, imag} */,
  {32'hc215830e, 32'h422b2d44} /* (22, 24, 23) {real, imag} */,
  {32'h42496623, 32'hc177631c} /* (22, 24, 22) {real, imag} */,
  {32'h42a13a3a, 32'h41a92c68} /* (22, 24, 21) {real, imag} */,
  {32'hc294ac79, 32'hc2815b64} /* (22, 24, 20) {real, imag} */,
  {32'hc2ffc44b, 32'hc2585584} /* (22, 24, 19) {real, imag} */,
  {32'hc0a4a69c, 32'h419833e3} /* (22, 24, 18) {real, imag} */,
  {32'h4236a799, 32'h42a677e2} /* (22, 24, 17) {real, imag} */,
  {32'hc2b387b2, 32'h00000000} /* (22, 24, 16) {real, imag} */,
  {32'h4236a799, 32'hc2a677e2} /* (22, 24, 15) {real, imag} */,
  {32'hc0a4a69c, 32'hc19833e3} /* (22, 24, 14) {real, imag} */,
  {32'hc2ffc44b, 32'h42585584} /* (22, 24, 13) {real, imag} */,
  {32'hc294ac79, 32'h42815b64} /* (22, 24, 12) {real, imag} */,
  {32'h42a13a3a, 32'hc1a92c68} /* (22, 24, 11) {real, imag} */,
  {32'h42496623, 32'h4177631c} /* (22, 24, 10) {real, imag} */,
  {32'hc215830e, 32'hc22b2d44} /* (22, 24, 9) {real, imag} */,
  {32'h428bacf6, 32'h423ae646} /* (22, 24, 8) {real, imag} */,
  {32'h423bc214, 32'hc2bbdd4e} /* (22, 24, 7) {real, imag} */,
  {32'h423f7984, 32'h420c71c7} /* (22, 24, 6) {real, imag} */,
  {32'h43501d60, 32'h4300e333} /* (22, 24, 5) {real, imag} */,
  {32'hc22e04c8, 32'hc3264515} /* (22, 24, 4) {real, imag} */,
  {32'hc2f992da, 32'hc28ca6b5} /* (22, 24, 3) {real, imag} */,
  {32'h44dd1d48, 32'h43428386} /* (22, 24, 2) {real, imag} */,
  {32'hc5848d57, 32'hc40c892a} /* (22, 24, 1) {real, imag} */,
  {32'hc5838923, 32'h00000000} /* (22, 24, 0) {real, imag} */,
  {32'hc55ac0c8, 32'h43cf228a} /* (22, 23, 31) {real, imag} */,
  {32'h44a6e68d, 32'hc3966fd9} /* (22, 23, 30) {real, imag} */,
  {32'h421dae5f, 32'hc2038af2} /* (22, 23, 29) {real, imag} */,
  {32'hc2a6284e, 32'h4329972b} /* (22, 23, 28) {real, imag} */,
  {32'h438065dc, 32'hc2a2ccc6} /* (22, 23, 27) {real, imag} */,
  {32'h41fc17ae, 32'hc30c4a24} /* (22, 23, 26) {real, imag} */,
  {32'h4198c467, 32'h427a2e46} /* (22, 23, 25) {real, imag} */,
  {32'h425b1c22, 32'h427d802c} /* (22, 23, 24) {real, imag} */,
  {32'hc23b0847, 32'hc234ad73} /* (22, 23, 23) {real, imag} */,
  {32'hc23204c9, 32'hc27f9fd0} /* (22, 23, 22) {real, imag} */,
  {32'hc05c8f28, 32'h4202dfdf} /* (22, 23, 21) {real, imag} */,
  {32'h41aab9b4, 32'h417b61ec} /* (22, 23, 20) {real, imag} */,
  {32'hc288ea0f, 32'hc28da21c} /* (22, 23, 19) {real, imag} */,
  {32'hc2292720, 32'h411f2a74} /* (22, 23, 18) {real, imag} */,
  {32'h4153f5aa, 32'hc1b85596} /* (22, 23, 17) {real, imag} */,
  {32'h427ff021, 32'h00000000} /* (22, 23, 16) {real, imag} */,
  {32'h4153f5aa, 32'h41b85596} /* (22, 23, 15) {real, imag} */,
  {32'hc2292720, 32'hc11f2a74} /* (22, 23, 14) {real, imag} */,
  {32'hc288ea0f, 32'h428da21c} /* (22, 23, 13) {real, imag} */,
  {32'h41aab9b4, 32'hc17b61ec} /* (22, 23, 12) {real, imag} */,
  {32'hc05c8f28, 32'hc202dfdf} /* (22, 23, 11) {real, imag} */,
  {32'hc23204c9, 32'h427f9fd0} /* (22, 23, 10) {real, imag} */,
  {32'hc23b0847, 32'h4234ad73} /* (22, 23, 9) {real, imag} */,
  {32'h425b1c22, 32'hc27d802c} /* (22, 23, 8) {real, imag} */,
  {32'h4198c467, 32'hc27a2e46} /* (22, 23, 7) {real, imag} */,
  {32'h41fc17ae, 32'h430c4a24} /* (22, 23, 6) {real, imag} */,
  {32'h438065dc, 32'h42a2ccc6} /* (22, 23, 5) {real, imag} */,
  {32'hc2a6284e, 32'hc329972b} /* (22, 23, 4) {real, imag} */,
  {32'h421dae5f, 32'h42038af2} /* (22, 23, 3) {real, imag} */,
  {32'h44a6e68d, 32'h43966fd9} /* (22, 23, 2) {real, imag} */,
  {32'hc55ac0c8, 32'hc3cf228a} /* (22, 23, 1) {real, imag} */,
  {32'hc55e7834, 32'h00000000} /* (22, 23, 0) {real, imag} */,
  {32'hc5177fbf, 32'h438eacca} /* (22, 22, 31) {real, imag} */,
  {32'h445734c4, 32'hc350bd50} /* (22, 22, 30) {real, imag} */,
  {32'h4197b3de, 32'h428e6952} /* (22, 22, 29) {real, imag} */,
  {32'hc30195f7, 32'h43374e45} /* (22, 22, 28) {real, imag} */,
  {32'h435019b9, 32'hc2ca67ae} /* (22, 22, 27) {real, imag} */,
  {32'hc118fea9, 32'hc2a418b2} /* (22, 22, 26) {real, imag} */,
  {32'hc2ae1bcc, 32'hc20ed82e} /* (22, 22, 25) {real, imag} */,
  {32'h42a50014, 32'hc253c684} /* (22, 22, 24) {real, imag} */,
  {32'h41b423d0, 32'h41210f62} /* (22, 22, 23) {real, imag} */,
  {32'hc240141d, 32'h41a1727b} /* (22, 22, 22) {real, imag} */,
  {32'h417fab36, 32'hc2afb028} /* (22, 22, 21) {real, imag} */,
  {32'h41b20219, 32'hc2bc7a6b} /* (22, 22, 20) {real, imag} */,
  {32'h41c7db74, 32'hc191101b} /* (22, 22, 19) {real, imag} */,
  {32'hc1d73348, 32'hc27b6f85} /* (22, 22, 18) {real, imag} */,
  {32'hc1a371d0, 32'h419e9491} /* (22, 22, 17) {real, imag} */,
  {32'h42796f0b, 32'h00000000} /* (22, 22, 16) {real, imag} */,
  {32'hc1a371d0, 32'hc19e9491} /* (22, 22, 15) {real, imag} */,
  {32'hc1d73348, 32'h427b6f85} /* (22, 22, 14) {real, imag} */,
  {32'h41c7db74, 32'h4191101b} /* (22, 22, 13) {real, imag} */,
  {32'h41b20219, 32'h42bc7a6b} /* (22, 22, 12) {real, imag} */,
  {32'h417fab36, 32'h42afb028} /* (22, 22, 11) {real, imag} */,
  {32'hc240141d, 32'hc1a1727b} /* (22, 22, 10) {real, imag} */,
  {32'h41b423d0, 32'hc1210f62} /* (22, 22, 9) {real, imag} */,
  {32'h42a50014, 32'h4253c684} /* (22, 22, 8) {real, imag} */,
  {32'hc2ae1bcc, 32'h420ed82e} /* (22, 22, 7) {real, imag} */,
  {32'hc118fea9, 32'h42a418b2} /* (22, 22, 6) {real, imag} */,
  {32'h435019b9, 32'h42ca67ae} /* (22, 22, 5) {real, imag} */,
  {32'hc30195f7, 32'hc3374e45} /* (22, 22, 4) {real, imag} */,
  {32'h4197b3de, 32'hc28e6952} /* (22, 22, 3) {real, imag} */,
  {32'h445734c4, 32'h4350bd50} /* (22, 22, 2) {real, imag} */,
  {32'hc5177fbf, 32'hc38eacca} /* (22, 22, 1) {real, imag} */,
  {32'hc51a84e4, 32'h00000000} /* (22, 22, 0) {real, imag} */,
  {32'hc46c99e0, 32'h42c373e4} /* (22, 21, 31) {real, imag} */,
  {32'h43896fd2, 32'hc33db3ef} /* (22, 21, 30) {real, imag} */,
  {32'h41feee68, 32'h431f189d} /* (22, 21, 29) {real, imag} */,
  {32'hc30bd2d9, 32'h42448b41} /* (22, 21, 28) {real, imag} */,
  {32'h4319cabf, 32'hc29299cc} /* (22, 21, 27) {real, imag} */,
  {32'hc2764f36, 32'h4105e1be} /* (22, 21, 26) {real, imag} */,
  {32'hc180c700, 32'hc2a84c92} /* (22, 21, 25) {real, imag} */,
  {32'h42f79728, 32'hc27c182b} /* (22, 21, 24) {real, imag} */,
  {32'hc2d80930, 32'h4214a110} /* (22, 21, 23) {real, imag} */,
  {32'h425068e8, 32'hc2993e68} /* (22, 21, 22) {real, imag} */,
  {32'h42648517, 32'hc24d6c45} /* (22, 21, 21) {real, imag} */,
  {32'h4186b200, 32'h42ae0060} /* (22, 21, 20) {real, imag} */,
  {32'h424b35b7, 32'hc24a81a7} /* (22, 21, 19) {real, imag} */,
  {32'hc2630931, 32'hc210aecc} /* (22, 21, 18) {real, imag} */,
  {32'h420ff327, 32'h423bdbdb} /* (22, 21, 17) {real, imag} */,
  {32'hc176afdb, 32'h00000000} /* (22, 21, 16) {real, imag} */,
  {32'h420ff327, 32'hc23bdbdb} /* (22, 21, 15) {real, imag} */,
  {32'hc2630931, 32'h4210aecc} /* (22, 21, 14) {real, imag} */,
  {32'h424b35b7, 32'h424a81a7} /* (22, 21, 13) {real, imag} */,
  {32'h4186b200, 32'hc2ae0060} /* (22, 21, 12) {real, imag} */,
  {32'h42648517, 32'h424d6c45} /* (22, 21, 11) {real, imag} */,
  {32'h425068e8, 32'h42993e68} /* (22, 21, 10) {real, imag} */,
  {32'hc2d80930, 32'hc214a110} /* (22, 21, 9) {real, imag} */,
  {32'h42f79728, 32'h427c182b} /* (22, 21, 8) {real, imag} */,
  {32'hc180c700, 32'h42a84c92} /* (22, 21, 7) {real, imag} */,
  {32'hc2764f36, 32'hc105e1be} /* (22, 21, 6) {real, imag} */,
  {32'h4319cabf, 32'h429299cc} /* (22, 21, 5) {real, imag} */,
  {32'hc30bd2d9, 32'hc2448b41} /* (22, 21, 4) {real, imag} */,
  {32'h41feee68, 32'hc31f189d} /* (22, 21, 3) {real, imag} */,
  {32'h43896fd2, 32'h433db3ef} /* (22, 21, 2) {real, imag} */,
  {32'hc46c99e0, 32'hc2c373e4} /* (22, 21, 1) {real, imag} */,
  {32'hc48e074e, 32'h00000000} /* (22, 21, 0) {real, imag} */,
  {32'h4491d7c4, 32'hc345bf4c} /* (22, 20, 31) {real, imag} */,
  {32'hc40f2b29, 32'hc2ca2ef5} /* (22, 20, 30) {real, imag} */,
  {32'hc29ecd36, 32'h42f4d36e} /* (22, 20, 29) {real, imag} */,
  {32'hc12b5ac0, 32'hc3076504} /* (22, 20, 28) {real, imag} */,
  {32'hc2dc4fd4, 32'hc1312f08} /* (22, 20, 27) {real, imag} */,
  {32'hc28e65b4, 32'hc3072828} /* (22, 20, 26) {real, imag} */,
  {32'h410ee10c, 32'h42738417} /* (22, 20, 25) {real, imag} */,
  {32'hc20cdcc3, 32'hc12b71c8} /* (22, 20, 24) {real, imag} */,
  {32'hc251afbe, 32'h4067f050} /* (22, 20, 23) {real, imag} */,
  {32'hc28fc8bf, 32'hc21d5aca} /* (22, 20, 22) {real, imag} */,
  {32'h41e270da, 32'h429c673c} /* (22, 20, 21) {real, imag} */,
  {32'h40efd668, 32'h42255a4e} /* (22, 20, 20) {real, imag} */,
  {32'h40114e94, 32'hc29f45fe} /* (22, 20, 19) {real, imag} */,
  {32'h416b4c2c, 32'h4193b7f0} /* (22, 20, 18) {real, imag} */,
  {32'h40248bb0, 32'h415aa362} /* (22, 20, 17) {real, imag} */,
  {32'h3f8d8d20, 32'h00000000} /* (22, 20, 16) {real, imag} */,
  {32'h40248bb0, 32'hc15aa362} /* (22, 20, 15) {real, imag} */,
  {32'h416b4c2c, 32'hc193b7f0} /* (22, 20, 14) {real, imag} */,
  {32'h40114e94, 32'h429f45fe} /* (22, 20, 13) {real, imag} */,
  {32'h40efd668, 32'hc2255a4e} /* (22, 20, 12) {real, imag} */,
  {32'h41e270da, 32'hc29c673c} /* (22, 20, 11) {real, imag} */,
  {32'hc28fc8bf, 32'h421d5aca} /* (22, 20, 10) {real, imag} */,
  {32'hc251afbe, 32'hc067f050} /* (22, 20, 9) {real, imag} */,
  {32'hc20cdcc3, 32'h412b71c8} /* (22, 20, 8) {real, imag} */,
  {32'h410ee10c, 32'hc2738417} /* (22, 20, 7) {real, imag} */,
  {32'hc28e65b4, 32'h43072828} /* (22, 20, 6) {real, imag} */,
  {32'hc2dc4fd4, 32'h41312f08} /* (22, 20, 5) {real, imag} */,
  {32'hc12b5ac0, 32'h43076504} /* (22, 20, 4) {real, imag} */,
  {32'hc29ecd36, 32'hc2f4d36e} /* (22, 20, 3) {real, imag} */,
  {32'hc40f2b29, 32'h42ca2ef5} /* (22, 20, 2) {real, imag} */,
  {32'h4491d7c4, 32'h4345bf4c} /* (22, 20, 1) {real, imag} */,
  {32'h43ea602c, 32'h00000000} /* (22, 20, 0) {real, imag} */,
  {32'h451a822a, 32'hc3be9b41} /* (22, 19, 31) {real, imag} */,
  {32'hc482e57e, 32'h43938af9} /* (22, 19, 30) {real, imag} */,
  {32'hc306263a, 32'h4264a838} /* (22, 19, 29) {real, imag} */,
  {32'h42b82e0c, 32'hc29aa04c} /* (22, 19, 28) {real, imag} */,
  {32'hc33d3235, 32'h4260f14c} /* (22, 19, 27) {real, imag} */,
  {32'h425f4b0d, 32'hc237d8e5} /* (22, 19, 26) {real, imag} */,
  {32'h4304613f, 32'h411c3858} /* (22, 19, 25) {real, imag} */,
  {32'hc2c26f76, 32'hc2cbddd8} /* (22, 19, 24) {real, imag} */,
  {32'h4235c4bb, 32'hc2806069} /* (22, 19, 23) {real, imag} */,
  {32'hc141e782, 32'h41815699} /* (22, 19, 22) {real, imag} */,
  {32'hc1218631, 32'h41883441} /* (22, 19, 21) {real, imag} */,
  {32'h41901da0, 32'h42409e0b} /* (22, 19, 20) {real, imag} */,
  {32'h4208641d, 32'hc2199c97} /* (22, 19, 19) {real, imag} */,
  {32'hc0c7f0e8, 32'hc23765e2} /* (22, 19, 18) {real, imag} */,
  {32'hbffb5fb8, 32'hc0f00bf4} /* (22, 19, 17) {real, imag} */,
  {32'hc28a1ff9, 32'h00000000} /* (22, 19, 16) {real, imag} */,
  {32'hbffb5fb8, 32'h40f00bf4} /* (22, 19, 15) {real, imag} */,
  {32'hc0c7f0e8, 32'h423765e2} /* (22, 19, 14) {real, imag} */,
  {32'h4208641d, 32'h42199c97} /* (22, 19, 13) {real, imag} */,
  {32'h41901da0, 32'hc2409e0b} /* (22, 19, 12) {real, imag} */,
  {32'hc1218631, 32'hc1883441} /* (22, 19, 11) {real, imag} */,
  {32'hc141e782, 32'hc1815699} /* (22, 19, 10) {real, imag} */,
  {32'h4235c4bb, 32'h42806069} /* (22, 19, 9) {real, imag} */,
  {32'hc2c26f76, 32'h42cbddd8} /* (22, 19, 8) {real, imag} */,
  {32'h4304613f, 32'hc11c3858} /* (22, 19, 7) {real, imag} */,
  {32'h425f4b0d, 32'h4237d8e5} /* (22, 19, 6) {real, imag} */,
  {32'hc33d3235, 32'hc260f14c} /* (22, 19, 5) {real, imag} */,
  {32'h42b82e0c, 32'h429aa04c} /* (22, 19, 4) {real, imag} */,
  {32'hc306263a, 32'hc264a838} /* (22, 19, 3) {real, imag} */,
  {32'hc482e57e, 32'hc3938af9} /* (22, 19, 2) {real, imag} */,
  {32'h451a822a, 32'h43be9b41} /* (22, 19, 1) {real, imag} */,
  {32'h44a335ac, 32'h00000000} /* (22, 19, 0) {real, imag} */,
  {32'h45588703, 32'hc3d48f9a} /* (22, 18, 31) {real, imag} */,
  {32'hc49f070b, 32'h439d94c8} /* (22, 18, 30) {real, imag} */,
  {32'hc2845c88, 32'hc2973c94} /* (22, 18, 29) {real, imag} */,
  {32'h4380142c, 32'hc307969e} /* (22, 18, 28) {real, imag} */,
  {32'hc21029aa, 32'h4330347c} /* (22, 18, 27) {real, imag} */,
  {32'hc2ae5c5d, 32'h4204155e} /* (22, 18, 26) {real, imag} */,
  {32'hc1c8d3d2, 32'hc23dffee} /* (22, 18, 25) {real, imag} */,
  {32'hbf376280, 32'h428b29d7} /* (22, 18, 24) {real, imag} */,
  {32'hc26ad8df, 32'hc1ec3521} /* (22, 18, 23) {real, imag} */,
  {32'hc1d11234, 32'h410eca1c} /* (22, 18, 22) {real, imag} */,
  {32'hc2581f18, 32'h4028a1c4} /* (22, 18, 21) {real, imag} */,
  {32'hc29132b8, 32'h423a4dc9} /* (22, 18, 20) {real, imag} */,
  {32'hc1ce8e07, 32'hc1ca9110} /* (22, 18, 19) {real, imag} */,
  {32'hc1988602, 32'h41f08e16} /* (22, 18, 18) {real, imag} */,
  {32'h425c2992, 32'h411888d5} /* (22, 18, 17) {real, imag} */,
  {32'hc17bd686, 32'h00000000} /* (22, 18, 16) {real, imag} */,
  {32'h425c2992, 32'hc11888d5} /* (22, 18, 15) {real, imag} */,
  {32'hc1988602, 32'hc1f08e16} /* (22, 18, 14) {real, imag} */,
  {32'hc1ce8e07, 32'h41ca9110} /* (22, 18, 13) {real, imag} */,
  {32'hc29132b8, 32'hc23a4dc9} /* (22, 18, 12) {real, imag} */,
  {32'hc2581f18, 32'hc028a1c4} /* (22, 18, 11) {real, imag} */,
  {32'hc1d11234, 32'hc10eca1c} /* (22, 18, 10) {real, imag} */,
  {32'hc26ad8df, 32'h41ec3521} /* (22, 18, 9) {real, imag} */,
  {32'hbf376280, 32'hc28b29d7} /* (22, 18, 8) {real, imag} */,
  {32'hc1c8d3d2, 32'h423dffee} /* (22, 18, 7) {real, imag} */,
  {32'hc2ae5c5d, 32'hc204155e} /* (22, 18, 6) {real, imag} */,
  {32'hc21029aa, 32'hc330347c} /* (22, 18, 5) {real, imag} */,
  {32'h4380142c, 32'h4307969e} /* (22, 18, 4) {real, imag} */,
  {32'hc2845c88, 32'h42973c94} /* (22, 18, 3) {real, imag} */,
  {32'hc49f070b, 32'hc39d94c8} /* (22, 18, 2) {real, imag} */,
  {32'h45588703, 32'h43d48f9a} /* (22, 18, 1) {real, imag} */,
  {32'h44f3bb48, 32'h00000000} /* (22, 18, 0) {real, imag} */,
  {32'h457e681b, 32'hc3cc9794} /* (22, 17, 31) {real, imag} */,
  {32'hc4bb3a38, 32'h43bcb830} /* (22, 17, 30) {real, imag} */,
  {32'hc1629f20, 32'h42895059} /* (22, 17, 29) {real, imag} */,
  {32'h43e31cd0, 32'hc3543ba0} /* (22, 17, 28) {real, imag} */,
  {32'hc3825f20, 32'h430ae443} /* (22, 17, 27) {real, imag} */,
  {32'hc29f2018, 32'hc22dea1c} /* (22, 17, 26) {real, imag} */,
  {32'h41d13d78, 32'h4277203e} /* (22, 17, 25) {real, imag} */,
  {32'h429a3f16, 32'h42dd19e9} /* (22, 17, 24) {real, imag} */,
  {32'hc192f442, 32'hc22a47f3} /* (22, 17, 23) {real, imag} */,
  {32'hc09bf602, 32'h429d6906} /* (22, 17, 22) {real, imag} */,
  {32'hc20083f2, 32'hc2aeeed1} /* (22, 17, 21) {real, imag} */,
  {32'hc25a2868, 32'h3fbf0340} /* (22, 17, 20) {real, imag} */,
  {32'hc21651ed, 32'h404bcaf0} /* (22, 17, 19) {real, imag} */,
  {32'hbf5b1700, 32'hc2b0cea1} /* (22, 17, 18) {real, imag} */,
  {32'h425b257e, 32'h4127afe6} /* (22, 17, 17) {real, imag} */,
  {32'hc18ef04e, 32'h00000000} /* (22, 17, 16) {real, imag} */,
  {32'h425b257e, 32'hc127afe6} /* (22, 17, 15) {real, imag} */,
  {32'hbf5b1700, 32'h42b0cea1} /* (22, 17, 14) {real, imag} */,
  {32'hc21651ed, 32'hc04bcaf0} /* (22, 17, 13) {real, imag} */,
  {32'hc25a2868, 32'hbfbf0340} /* (22, 17, 12) {real, imag} */,
  {32'hc20083f2, 32'h42aeeed1} /* (22, 17, 11) {real, imag} */,
  {32'hc09bf602, 32'hc29d6906} /* (22, 17, 10) {real, imag} */,
  {32'hc192f442, 32'h422a47f3} /* (22, 17, 9) {real, imag} */,
  {32'h429a3f16, 32'hc2dd19e9} /* (22, 17, 8) {real, imag} */,
  {32'h41d13d78, 32'hc277203e} /* (22, 17, 7) {real, imag} */,
  {32'hc29f2018, 32'h422dea1c} /* (22, 17, 6) {real, imag} */,
  {32'hc3825f20, 32'hc30ae443} /* (22, 17, 5) {real, imag} */,
  {32'h43e31cd0, 32'h43543ba0} /* (22, 17, 4) {real, imag} */,
  {32'hc1629f20, 32'hc2895059} /* (22, 17, 3) {real, imag} */,
  {32'hc4bb3a38, 32'hc3bcb830} /* (22, 17, 2) {real, imag} */,
  {32'h457e681b, 32'h43cc9794} /* (22, 17, 1) {real, imag} */,
  {32'h451eee1c, 32'h00000000} /* (22, 17, 0) {real, imag} */,
  {32'h4585459a, 32'hc3df07ac} /* (22, 16, 31) {real, imag} */,
  {32'hc4bf009f, 32'h438e3925} /* (22, 16, 30) {real, imag} */,
  {32'hc29feb8a, 32'h437211a0} /* (22, 16, 29) {real, imag} */,
  {32'h43ccfc3c, 32'hc38e6fc8} /* (22, 16, 28) {real, imag} */,
  {32'hc3848297, 32'h4292aae2} /* (22, 16, 27) {real, imag} */,
  {32'hc27508e4, 32'hc2a42723} /* (22, 16, 26) {real, imag} */,
  {32'h425901bf, 32'hc25f649a} /* (22, 16, 25) {real, imag} */,
  {32'hc26ffaa8, 32'h4257deec} /* (22, 16, 24) {real, imag} */,
  {32'hc21528b6, 32'h414e8f50} /* (22, 16, 23) {real, imag} */,
  {32'h42c77f0d, 32'h41555a54} /* (22, 16, 22) {real, imag} */,
  {32'h41a2ebd4, 32'hc203a66d} /* (22, 16, 21) {real, imag} */,
  {32'hc29f4127, 32'h4321e6de} /* (22, 16, 20) {real, imag} */,
  {32'hc19e19c4, 32'hc1fd21a0} /* (22, 16, 19) {real, imag} */,
  {32'h403c47d8, 32'h42239db5} /* (22, 16, 18) {real, imag} */,
  {32'hc1b8f861, 32'hc1277320} /* (22, 16, 17) {real, imag} */,
  {32'hc24c7e3f, 32'h00000000} /* (22, 16, 16) {real, imag} */,
  {32'hc1b8f861, 32'h41277320} /* (22, 16, 15) {real, imag} */,
  {32'h403c47d8, 32'hc2239db5} /* (22, 16, 14) {real, imag} */,
  {32'hc19e19c4, 32'h41fd21a0} /* (22, 16, 13) {real, imag} */,
  {32'hc29f4127, 32'hc321e6de} /* (22, 16, 12) {real, imag} */,
  {32'h41a2ebd4, 32'h4203a66d} /* (22, 16, 11) {real, imag} */,
  {32'h42c77f0d, 32'hc1555a54} /* (22, 16, 10) {real, imag} */,
  {32'hc21528b6, 32'hc14e8f50} /* (22, 16, 9) {real, imag} */,
  {32'hc26ffaa8, 32'hc257deec} /* (22, 16, 8) {real, imag} */,
  {32'h425901bf, 32'h425f649a} /* (22, 16, 7) {real, imag} */,
  {32'hc27508e4, 32'h42a42723} /* (22, 16, 6) {real, imag} */,
  {32'hc3848297, 32'hc292aae2} /* (22, 16, 5) {real, imag} */,
  {32'h43ccfc3c, 32'h438e6fc8} /* (22, 16, 4) {real, imag} */,
  {32'hc29feb8a, 32'hc37211a0} /* (22, 16, 3) {real, imag} */,
  {32'hc4bf009f, 32'hc38e3925} /* (22, 16, 2) {real, imag} */,
  {32'h4585459a, 32'h43df07ac} /* (22, 16, 1) {real, imag} */,
  {32'h452e8e02, 32'h00000000} /* (22, 16, 0) {real, imag} */,
  {32'h4585a3e2, 32'hc3bc6b64} /* (22, 15, 31) {real, imag} */,
  {32'hc4b37df4, 32'h43965eec} /* (22, 15, 30) {real, imag} */,
  {32'hc35fdf80, 32'h430c902e} /* (22, 15, 29) {real, imag} */,
  {32'h43949784, 32'hc3588df6} /* (22, 15, 28) {real, imag} */,
  {32'hc386155e, 32'h43237639} /* (22, 15, 27) {real, imag} */,
  {32'hc359468c, 32'hc192702c} /* (22, 15, 26) {real, imag} */,
  {32'h42d48c7a, 32'hc29af241} /* (22, 15, 25) {real, imag} */,
  {32'hc1c46bd6, 32'h425a84f6} /* (22, 15, 24) {real, imag} */,
  {32'h411d40db, 32'h400785b0} /* (22, 15, 23) {real, imag} */,
  {32'hc11d0301, 32'hc15e68d0} /* (22, 15, 22) {real, imag} */,
  {32'hbfde4638, 32'h42caffdf} /* (22, 15, 21) {real, imag} */,
  {32'hc1f07297, 32'hc2096012} /* (22, 15, 20) {real, imag} */,
  {32'h4127b4b5, 32'h42924a64} /* (22, 15, 19) {real, imag} */,
  {32'hc22f5846, 32'h406e3020} /* (22, 15, 18) {real, imag} */,
  {32'h3db92900, 32'h408e1011} /* (22, 15, 17) {real, imag} */,
  {32'h41c69d24, 32'h00000000} /* (22, 15, 16) {real, imag} */,
  {32'h3db92900, 32'hc08e1011} /* (22, 15, 15) {real, imag} */,
  {32'hc22f5846, 32'hc06e3020} /* (22, 15, 14) {real, imag} */,
  {32'h4127b4b5, 32'hc2924a64} /* (22, 15, 13) {real, imag} */,
  {32'hc1f07297, 32'h42096012} /* (22, 15, 12) {real, imag} */,
  {32'hbfde4638, 32'hc2caffdf} /* (22, 15, 11) {real, imag} */,
  {32'hc11d0301, 32'h415e68d0} /* (22, 15, 10) {real, imag} */,
  {32'h411d40db, 32'hc00785b0} /* (22, 15, 9) {real, imag} */,
  {32'hc1c46bd6, 32'hc25a84f6} /* (22, 15, 8) {real, imag} */,
  {32'h42d48c7a, 32'h429af241} /* (22, 15, 7) {real, imag} */,
  {32'hc359468c, 32'h4192702c} /* (22, 15, 6) {real, imag} */,
  {32'hc386155e, 32'hc3237639} /* (22, 15, 5) {real, imag} */,
  {32'h43949784, 32'h43588df6} /* (22, 15, 4) {real, imag} */,
  {32'hc35fdf80, 32'hc30c902e} /* (22, 15, 3) {real, imag} */,
  {32'hc4b37df4, 32'hc3965eec} /* (22, 15, 2) {real, imag} */,
  {32'h4585a3e2, 32'h43bc6b64} /* (22, 15, 1) {real, imag} */,
  {32'h45332340, 32'h00000000} /* (22, 15, 0) {real, imag} */,
  {32'h457535e5, 32'hc3b214fe} /* (22, 14, 31) {real, imag} */,
  {32'hc4bb22f3, 32'h437af3b4} /* (22, 14, 30) {real, imag} */,
  {32'hc282fcce, 32'h424ba4ad} /* (22, 14, 29) {real, imag} */,
  {32'h43ca1be0, 32'hc30cce7a} /* (22, 14, 28) {real, imag} */,
  {32'hc352edf0, 32'h42ad9a28} /* (22, 14, 27) {real, imag} */,
  {32'hc2b5b4d7, 32'hc130fe20} /* (22, 14, 26) {real, imag} */,
  {32'h42fc3540, 32'hc25f2742} /* (22, 14, 25) {real, imag} */,
  {32'hc2eb611f, 32'h408d32d0} /* (22, 14, 24) {real, imag} */,
  {32'h4254ea1b, 32'h42b24681} /* (22, 14, 23) {real, imag} */,
  {32'h430a64a0, 32'h42fbb162} /* (22, 14, 22) {real, imag} */,
  {32'hc18e4317, 32'hc1a3428e} /* (22, 14, 21) {real, imag} */,
  {32'h414fe964, 32'h42a80758} /* (22, 14, 20) {real, imag} */,
  {32'h404612b8, 32'hc20144d7} /* (22, 14, 19) {real, imag} */,
  {32'h423d59fb, 32'h425f7fc9} /* (22, 14, 18) {real, imag} */,
  {32'h423a286c, 32'hc103804f} /* (22, 14, 17) {real, imag} */,
  {32'h421f13ee, 32'h00000000} /* (22, 14, 16) {real, imag} */,
  {32'h423a286c, 32'h4103804f} /* (22, 14, 15) {real, imag} */,
  {32'h423d59fb, 32'hc25f7fc9} /* (22, 14, 14) {real, imag} */,
  {32'h404612b8, 32'h420144d7} /* (22, 14, 13) {real, imag} */,
  {32'h414fe964, 32'hc2a80758} /* (22, 14, 12) {real, imag} */,
  {32'hc18e4317, 32'h41a3428e} /* (22, 14, 11) {real, imag} */,
  {32'h430a64a0, 32'hc2fbb162} /* (22, 14, 10) {real, imag} */,
  {32'h4254ea1b, 32'hc2b24681} /* (22, 14, 9) {real, imag} */,
  {32'hc2eb611f, 32'hc08d32d0} /* (22, 14, 8) {real, imag} */,
  {32'h42fc3540, 32'h425f2742} /* (22, 14, 7) {real, imag} */,
  {32'hc2b5b4d7, 32'h4130fe20} /* (22, 14, 6) {real, imag} */,
  {32'hc352edf0, 32'hc2ad9a28} /* (22, 14, 5) {real, imag} */,
  {32'h43ca1be0, 32'h430cce7a} /* (22, 14, 4) {real, imag} */,
  {32'hc282fcce, 32'hc24ba4ad} /* (22, 14, 3) {real, imag} */,
  {32'hc4bb22f3, 32'hc37af3b4} /* (22, 14, 2) {real, imag} */,
  {32'h457535e5, 32'h43b214fe} /* (22, 14, 1) {real, imag} */,
  {32'h45379dc4, 32'h00000000} /* (22, 14, 0) {real, imag} */,
  {32'h454f5b7c, 32'hbd61e000} /* (22, 13, 31) {real, imag} */,
  {32'hc4b24bbe, 32'h43113430} /* (22, 13, 30) {real, imag} */,
  {32'hc1d5bfce, 32'hc1e30ee8} /* (22, 13, 29) {real, imag} */,
  {32'h439ccdaf, 32'hc37bfd6e} /* (22, 13, 28) {real, imag} */,
  {32'hc33f1d3f, 32'h43641c5b} /* (22, 13, 27) {real, imag} */,
  {32'h401a4550, 32'hc27816cb} /* (22, 13, 26) {real, imag} */,
  {32'h42830034, 32'hc2ec17b9} /* (22, 13, 25) {real, imag} */,
  {32'hc2cec5b8, 32'h4322c8aa} /* (22, 13, 24) {real, imag} */,
  {32'h42549231, 32'h42931285} /* (22, 13, 23) {real, imag} */,
  {32'h42198dcc, 32'hc196586b} /* (22, 13, 22) {real, imag} */,
  {32'hc101c7fb, 32'h42152e54} /* (22, 13, 21) {real, imag} */,
  {32'hc238baa6, 32'hc192c62a} /* (22, 13, 20) {real, imag} */,
  {32'h4299fe02, 32'h419ba1e2} /* (22, 13, 19) {real, imag} */,
  {32'hc10ca0ac, 32'h42888e0f} /* (22, 13, 18) {real, imag} */,
  {32'hbfa3c488, 32'h421c2f54} /* (22, 13, 17) {real, imag} */,
  {32'h422d8bca, 32'h00000000} /* (22, 13, 16) {real, imag} */,
  {32'hbfa3c488, 32'hc21c2f54} /* (22, 13, 15) {real, imag} */,
  {32'hc10ca0ac, 32'hc2888e0f} /* (22, 13, 14) {real, imag} */,
  {32'h4299fe02, 32'hc19ba1e2} /* (22, 13, 13) {real, imag} */,
  {32'hc238baa6, 32'h4192c62a} /* (22, 13, 12) {real, imag} */,
  {32'hc101c7fb, 32'hc2152e54} /* (22, 13, 11) {real, imag} */,
  {32'h42198dcc, 32'h4196586b} /* (22, 13, 10) {real, imag} */,
  {32'h42549231, 32'hc2931285} /* (22, 13, 9) {real, imag} */,
  {32'hc2cec5b8, 32'hc322c8aa} /* (22, 13, 8) {real, imag} */,
  {32'h42830034, 32'h42ec17b9} /* (22, 13, 7) {real, imag} */,
  {32'h401a4550, 32'h427816cb} /* (22, 13, 6) {real, imag} */,
  {32'hc33f1d3f, 32'hc3641c5b} /* (22, 13, 5) {real, imag} */,
  {32'h439ccdaf, 32'h437bfd6e} /* (22, 13, 4) {real, imag} */,
  {32'hc1d5bfce, 32'h41e30ee8} /* (22, 13, 3) {real, imag} */,
  {32'hc4b24bbe, 32'hc3113430} /* (22, 13, 2) {real, imag} */,
  {32'h454f5b7c, 32'h3d61e000} /* (22, 13, 1) {real, imag} */,
  {32'h451e6b6e, 32'h00000000} /* (22, 13, 0) {real, imag} */,
  {32'h45174166, 32'h432a20fc} /* (22, 12, 31) {real, imag} */,
  {32'hc49de9e2, 32'h429464c5} /* (22, 12, 30) {real, imag} */,
  {32'hc2b82142, 32'h42cdfd56} /* (22, 12, 29) {real, imag} */,
  {32'h437ef67a, 32'hc3907bc6} /* (22, 12, 28) {real, imag} */,
  {32'hc397aac2, 32'h4329036e} /* (22, 12, 27) {real, imag} */,
  {32'h42eed624, 32'h42c48754} /* (22, 12, 26) {real, imag} */,
  {32'h42c30bce, 32'h41c7f6ea} /* (22, 12, 25) {real, imag} */,
  {32'hc2b5a86e, 32'h40269420} /* (22, 12, 24) {real, imag} */,
  {32'hc144de50, 32'hc2defcfe} /* (22, 12, 23) {real, imag} */,
  {32'hc25b3c23, 32'h4240bc3c} /* (22, 12, 22) {real, imag} */,
  {32'hc288ce3c, 32'hc21fc3d9} /* (22, 12, 21) {real, imag} */,
  {32'hc289676a, 32'hc2bd97b7} /* (22, 12, 20) {real, imag} */,
  {32'h4208c0b4, 32'h42d3846c} /* (22, 12, 19) {real, imag} */,
  {32'hc246f879, 32'h412b6d9b} /* (22, 12, 18) {real, imag} */,
  {32'hc22a7cbd, 32'h4061bb48} /* (22, 12, 17) {real, imag} */,
  {32'hc293d100, 32'h00000000} /* (22, 12, 16) {real, imag} */,
  {32'hc22a7cbd, 32'hc061bb48} /* (22, 12, 15) {real, imag} */,
  {32'hc246f879, 32'hc12b6d9b} /* (22, 12, 14) {real, imag} */,
  {32'h4208c0b4, 32'hc2d3846c} /* (22, 12, 13) {real, imag} */,
  {32'hc289676a, 32'h42bd97b7} /* (22, 12, 12) {real, imag} */,
  {32'hc288ce3c, 32'h421fc3d9} /* (22, 12, 11) {real, imag} */,
  {32'hc25b3c23, 32'hc240bc3c} /* (22, 12, 10) {real, imag} */,
  {32'hc144de50, 32'h42defcfe} /* (22, 12, 9) {real, imag} */,
  {32'hc2b5a86e, 32'hc0269420} /* (22, 12, 8) {real, imag} */,
  {32'h42c30bce, 32'hc1c7f6ea} /* (22, 12, 7) {real, imag} */,
  {32'h42eed624, 32'hc2c48754} /* (22, 12, 6) {real, imag} */,
  {32'hc397aac2, 32'hc329036e} /* (22, 12, 5) {real, imag} */,
  {32'h437ef67a, 32'h43907bc6} /* (22, 12, 4) {real, imag} */,
  {32'hc2b82142, 32'hc2cdfd56} /* (22, 12, 3) {real, imag} */,
  {32'hc49de9e2, 32'hc29464c5} /* (22, 12, 2) {real, imag} */,
  {32'h45174166, 32'hc32a20fc} /* (22, 12, 1) {real, imag} */,
  {32'h44d7b7e9, 32'h00000000} /* (22, 12, 0) {real, imag} */,
  {32'h4493a188, 32'h43e0f843} /* (22, 11, 31) {real, imag} */,
  {32'hc44bca6d, 32'h3e6e2c00} /* (22, 11, 30) {real, imag} */,
  {32'hc2be43f8, 32'h41b0bf08} /* (22, 11, 29) {real, imag} */,
  {32'h43a03258, 32'hc25b1e2d} /* (22, 11, 28) {real, imag} */,
  {32'hc311afb7, 32'h42ef338e} /* (22, 11, 27) {real, imag} */,
  {32'hc1d84e01, 32'h424c07aa} /* (22, 11, 26) {real, imag} */,
  {32'h42d60a3d, 32'hc2d7ab96} /* (22, 11, 25) {real, imag} */,
  {32'hc20e2b49, 32'hc2446b51} /* (22, 11, 24) {real, imag} */,
  {32'h4296219e, 32'h4280b86a} /* (22, 11, 23) {real, imag} */,
  {32'hc16815e0, 32'h42f71efa} /* (22, 11, 22) {real, imag} */,
  {32'hc27ea41b, 32'hc0864eb8} /* (22, 11, 21) {real, imag} */,
  {32'h42a22e0b, 32'hc2c500f4} /* (22, 11, 20) {real, imag} */,
  {32'h41a0694e, 32'h415c1aec} /* (22, 11, 19) {real, imag} */,
  {32'hc28093d8, 32'h42843e1c} /* (22, 11, 18) {real, imag} */,
  {32'hc13fbfb4, 32'h41892642} /* (22, 11, 17) {real, imag} */,
  {32'h4163b1e1, 32'h00000000} /* (22, 11, 16) {real, imag} */,
  {32'hc13fbfb4, 32'hc1892642} /* (22, 11, 15) {real, imag} */,
  {32'hc28093d8, 32'hc2843e1c} /* (22, 11, 14) {real, imag} */,
  {32'h41a0694e, 32'hc15c1aec} /* (22, 11, 13) {real, imag} */,
  {32'h42a22e0b, 32'h42c500f4} /* (22, 11, 12) {real, imag} */,
  {32'hc27ea41b, 32'h40864eb8} /* (22, 11, 11) {real, imag} */,
  {32'hc16815e0, 32'hc2f71efa} /* (22, 11, 10) {real, imag} */,
  {32'h4296219e, 32'hc280b86a} /* (22, 11, 9) {real, imag} */,
  {32'hc20e2b49, 32'h42446b51} /* (22, 11, 8) {real, imag} */,
  {32'h42d60a3d, 32'h42d7ab96} /* (22, 11, 7) {real, imag} */,
  {32'hc1d84e01, 32'hc24c07aa} /* (22, 11, 6) {real, imag} */,
  {32'hc311afb7, 32'hc2ef338e} /* (22, 11, 5) {real, imag} */,
  {32'h43a03258, 32'h425b1e2d} /* (22, 11, 4) {real, imag} */,
  {32'hc2be43f8, 32'hc1b0bf08} /* (22, 11, 3) {real, imag} */,
  {32'hc44bca6d, 32'hbe6e2c00} /* (22, 11, 2) {real, imag} */,
  {32'h4493a188, 32'hc3e0f843} /* (22, 11, 1) {real, imag} */,
  {32'h4410fdac, 32'h00000000} /* (22, 11, 0) {real, imag} */,
  {32'hc422cd29, 32'h444e4ca1} /* (22, 10, 31) {real, imag} */,
  {32'h42020f38, 32'hc32a2f4a} /* (22, 10, 30) {real, imag} */,
  {32'hc194993a, 32'hc25745de} /* (22, 10, 29) {real, imag} */,
  {32'h42c2892e, 32'h431c3181} /* (22, 10, 28) {real, imag} */,
  {32'h430c48af, 32'hbf8ea1e0} /* (22, 10, 27) {real, imag} */,
  {32'h420199d2, 32'h4294bd64} /* (22, 10, 26) {real, imag} */,
  {32'h41f8d75a, 32'h41549fda} /* (22, 10, 25) {real, imag} */,
  {32'h4228e334, 32'hc2ca73c2} /* (22, 10, 24) {real, imag} */,
  {32'hc192ef78, 32'h4283fe5c} /* (22, 10, 23) {real, imag} */,
  {32'h4279d0ab, 32'h423bc410} /* (22, 10, 22) {real, imag} */,
  {32'hc2452bae, 32'hc2a9a566} /* (22, 10, 21) {real, imag} */,
  {32'h41f56347, 32'h429df69d} /* (22, 10, 20) {real, imag} */,
  {32'h423ddd0a, 32'h40a9e8a4} /* (22, 10, 19) {real, imag} */,
  {32'hc297dc7f, 32'h41ed061e} /* (22, 10, 18) {real, imag} */,
  {32'hc1ecd81c, 32'h42320b6c} /* (22, 10, 17) {real, imag} */,
  {32'h41b5124a, 32'h00000000} /* (22, 10, 16) {real, imag} */,
  {32'hc1ecd81c, 32'hc2320b6c} /* (22, 10, 15) {real, imag} */,
  {32'hc297dc7f, 32'hc1ed061e} /* (22, 10, 14) {real, imag} */,
  {32'h423ddd0a, 32'hc0a9e8a4} /* (22, 10, 13) {real, imag} */,
  {32'h41f56347, 32'hc29df69d} /* (22, 10, 12) {real, imag} */,
  {32'hc2452bae, 32'h42a9a566} /* (22, 10, 11) {real, imag} */,
  {32'h4279d0ab, 32'hc23bc410} /* (22, 10, 10) {real, imag} */,
  {32'hc192ef78, 32'hc283fe5c} /* (22, 10, 9) {real, imag} */,
  {32'h4228e334, 32'h42ca73c2} /* (22, 10, 8) {real, imag} */,
  {32'h41f8d75a, 32'hc1549fda} /* (22, 10, 7) {real, imag} */,
  {32'h420199d2, 32'hc294bd64} /* (22, 10, 6) {real, imag} */,
  {32'h430c48af, 32'h3f8ea1e0} /* (22, 10, 5) {real, imag} */,
  {32'h42c2892e, 32'hc31c3181} /* (22, 10, 4) {real, imag} */,
  {32'hc194993a, 32'h425745de} /* (22, 10, 3) {real, imag} */,
  {32'h42020f38, 32'h432a2f4a} /* (22, 10, 2) {real, imag} */,
  {32'hc422cd29, 32'hc44e4ca1} /* (22, 10, 1) {real, imag} */,
  {32'hc4655a96, 32'h00000000} /* (22, 10, 0) {real, imag} */,
  {32'hc50a79b4, 32'h448a5f02} /* (22, 9, 31) {real, imag} */,
  {32'h4409ec0a, 32'hc3dd6491} /* (22, 9, 30) {real, imag} */,
  {32'hc22b697d, 32'hc1f3c9a8} /* (22, 9, 29) {real, imag} */,
  {32'h4131f444, 32'h430a3d75} /* (22, 9, 28) {real, imag} */,
  {32'h4309a9d6, 32'hc32bf506} /* (22, 9, 27) {real, imag} */,
  {32'h420f079b, 32'h41ef48e4} /* (22, 9, 26) {real, imag} */,
  {32'h3fd3da70, 32'h4183aadc} /* (22, 9, 25) {real, imag} */,
  {32'h41916e77, 32'hc12e7772} /* (22, 9, 24) {real, imag} */,
  {32'hc26523e3, 32'h41cfc89a} /* (22, 9, 23) {real, imag} */,
  {32'hc2378787, 32'hc2cb04da} /* (22, 9, 22) {real, imag} */,
  {32'hc27924b4, 32'hc2ef4fb6} /* (22, 9, 21) {real, imag} */,
  {32'h418316f0, 32'hc2d25d62} /* (22, 9, 20) {real, imag} */,
  {32'h41853b1f, 32'h4211f21b} /* (22, 9, 19) {real, imag} */,
  {32'h41aef6d0, 32'hc2ee20c6} /* (22, 9, 18) {real, imag} */,
  {32'h3f89d904, 32'h41830c62} /* (22, 9, 17) {real, imag} */,
  {32'h424ee867, 32'h00000000} /* (22, 9, 16) {real, imag} */,
  {32'h3f89d904, 32'hc1830c62} /* (22, 9, 15) {real, imag} */,
  {32'h41aef6d0, 32'h42ee20c6} /* (22, 9, 14) {real, imag} */,
  {32'h41853b1f, 32'hc211f21b} /* (22, 9, 13) {real, imag} */,
  {32'h418316f0, 32'h42d25d62} /* (22, 9, 12) {real, imag} */,
  {32'hc27924b4, 32'h42ef4fb6} /* (22, 9, 11) {real, imag} */,
  {32'hc2378787, 32'h42cb04da} /* (22, 9, 10) {real, imag} */,
  {32'hc26523e3, 32'hc1cfc89a} /* (22, 9, 9) {real, imag} */,
  {32'h41916e77, 32'h412e7772} /* (22, 9, 8) {real, imag} */,
  {32'h3fd3da70, 32'hc183aadc} /* (22, 9, 7) {real, imag} */,
  {32'h420f079b, 32'hc1ef48e4} /* (22, 9, 6) {real, imag} */,
  {32'h4309a9d6, 32'h432bf506} /* (22, 9, 5) {real, imag} */,
  {32'h4131f444, 32'hc30a3d75} /* (22, 9, 4) {real, imag} */,
  {32'hc22b697d, 32'h41f3c9a8} /* (22, 9, 3) {real, imag} */,
  {32'h4409ec0a, 32'h43dd6491} /* (22, 9, 2) {real, imag} */,
  {32'hc50a79b4, 32'hc48a5f02} /* (22, 9, 1) {real, imag} */,
  {32'hc50f16cc, 32'h00000000} /* (22, 9, 0) {real, imag} */,
  {32'hc53c90a8, 32'h44c0451d} /* (22, 8, 31) {real, imag} */,
  {32'h447b90c0, 32'hc3de17eb} /* (22, 8, 30) {real, imag} */,
  {32'h404b5e50, 32'hc2b671df} /* (22, 8, 29) {real, imag} */,
  {32'hc300afa6, 32'h42c18d66} /* (22, 8, 28) {real, imag} */,
  {32'h435b6dec, 32'hc228092c} /* (22, 8, 27) {real, imag} */,
  {32'h4280a381, 32'h41800b74} /* (22, 8, 26) {real, imag} */,
  {32'h428d2883, 32'hc1dd83e8} /* (22, 8, 25) {real, imag} */,
  {32'hc212ed6a, 32'hc23d62ca} /* (22, 8, 24) {real, imag} */,
  {32'h432d155e, 32'hc20d9aa0} /* (22, 8, 23) {real, imag} */,
  {32'h41b23d3a, 32'h410b7894} /* (22, 8, 22) {real, imag} */,
  {32'h4265130b, 32'hc2ce0b47} /* (22, 8, 21) {real, imag} */,
  {32'hc15893d6, 32'h42756c40} /* (22, 8, 20) {real, imag} */,
  {32'h42e3ff75, 32'h41cacf65} /* (22, 8, 19) {real, imag} */,
  {32'h420fc338, 32'h4175d9f2} /* (22, 8, 18) {real, imag} */,
  {32'hc23001a7, 32'hc0eca2e0} /* (22, 8, 17) {real, imag} */,
  {32'h40bd0d80, 32'h00000000} /* (22, 8, 16) {real, imag} */,
  {32'hc23001a7, 32'h40eca2e0} /* (22, 8, 15) {real, imag} */,
  {32'h420fc338, 32'hc175d9f2} /* (22, 8, 14) {real, imag} */,
  {32'h42e3ff75, 32'hc1cacf65} /* (22, 8, 13) {real, imag} */,
  {32'hc15893d6, 32'hc2756c40} /* (22, 8, 12) {real, imag} */,
  {32'h4265130b, 32'h42ce0b47} /* (22, 8, 11) {real, imag} */,
  {32'h41b23d3a, 32'hc10b7894} /* (22, 8, 10) {real, imag} */,
  {32'h432d155e, 32'h420d9aa0} /* (22, 8, 9) {real, imag} */,
  {32'hc212ed6a, 32'h423d62ca} /* (22, 8, 8) {real, imag} */,
  {32'h428d2883, 32'h41dd83e8} /* (22, 8, 7) {real, imag} */,
  {32'h4280a381, 32'hc1800b74} /* (22, 8, 6) {real, imag} */,
  {32'h435b6dec, 32'h4228092c} /* (22, 8, 5) {real, imag} */,
  {32'hc300afa6, 32'hc2c18d66} /* (22, 8, 4) {real, imag} */,
  {32'h404b5e50, 32'h42b671df} /* (22, 8, 3) {real, imag} */,
  {32'h447b90c0, 32'h43de17eb} /* (22, 8, 2) {real, imag} */,
  {32'hc53c90a8, 32'hc4c0451d} /* (22, 8, 1) {real, imag} */,
  {32'hc54d750e, 32'h00000000} /* (22, 8, 0) {real, imag} */,
  {32'hc55e4f94, 32'h44fa7ee8} /* (22, 7, 31) {real, imag} */,
  {32'h4476ef49, 32'hc40f5ad1} /* (22, 7, 30) {real, imag} */,
  {32'h42a49e49, 32'hc2f24126} /* (22, 7, 29) {real, imag} */,
  {32'hc29b4202, 32'h426aa824} /* (22, 7, 28) {real, imag} */,
  {32'h4361f3b1, 32'hc1a5ce06} /* (22, 7, 27) {real, imag} */,
  {32'h40c77848, 32'h420c9220} /* (22, 7, 26) {real, imag} */,
  {32'h42b1029b, 32'hc24802f6} /* (22, 7, 25) {real, imag} */,
  {32'h42c0651d, 32'hc2e0589c} /* (22, 7, 24) {real, imag} */,
  {32'h41f1b2da, 32'hc24f70de} /* (22, 7, 23) {real, imag} */,
  {32'h427874ad, 32'h42fc4cd1} /* (22, 7, 22) {real, imag} */,
  {32'h428b93e0, 32'h41f8a262} /* (22, 7, 21) {real, imag} */,
  {32'hc2359623, 32'h42a4e6c4} /* (22, 7, 20) {real, imag} */,
  {32'hc2b4a979, 32'hc2aa1128} /* (22, 7, 19) {real, imag} */,
  {32'hc2cbe024, 32'hc2629c28} /* (22, 7, 18) {real, imag} */,
  {32'h41a6bbd4, 32'h41790e09} /* (22, 7, 17) {real, imag} */,
  {32'hc1b5f9cb, 32'h00000000} /* (22, 7, 16) {real, imag} */,
  {32'h41a6bbd4, 32'hc1790e09} /* (22, 7, 15) {real, imag} */,
  {32'hc2cbe024, 32'h42629c28} /* (22, 7, 14) {real, imag} */,
  {32'hc2b4a979, 32'h42aa1128} /* (22, 7, 13) {real, imag} */,
  {32'hc2359623, 32'hc2a4e6c4} /* (22, 7, 12) {real, imag} */,
  {32'h428b93e0, 32'hc1f8a262} /* (22, 7, 11) {real, imag} */,
  {32'h427874ad, 32'hc2fc4cd1} /* (22, 7, 10) {real, imag} */,
  {32'h41f1b2da, 32'h424f70de} /* (22, 7, 9) {real, imag} */,
  {32'h42c0651d, 32'h42e0589c} /* (22, 7, 8) {real, imag} */,
  {32'h42b1029b, 32'h424802f6} /* (22, 7, 7) {real, imag} */,
  {32'h40c77848, 32'hc20c9220} /* (22, 7, 6) {real, imag} */,
  {32'h4361f3b1, 32'h41a5ce06} /* (22, 7, 5) {real, imag} */,
  {32'hc29b4202, 32'hc26aa824} /* (22, 7, 4) {real, imag} */,
  {32'h42a49e49, 32'h42f24126} /* (22, 7, 3) {real, imag} */,
  {32'h4476ef49, 32'h440f5ad1} /* (22, 7, 2) {real, imag} */,
  {32'hc55e4f94, 32'hc4fa7ee8} /* (22, 7, 1) {real, imag} */,
  {32'hc57dfa91, 32'h00000000} /* (22, 7, 0) {real, imag} */,
  {32'hc5690f08, 32'h451c4712} /* (22, 6, 31) {real, imag} */,
  {32'h44476cb4, 32'hc4184eec} /* (22, 6, 30) {real, imag} */,
  {32'h428e0fea, 32'hc155220c} /* (22, 6, 29) {real, imag} */,
  {32'hc2437b90, 32'hc2a04fae} /* (22, 6, 28) {real, imag} */,
  {32'h43041655, 32'hc29f6f6f} /* (22, 6, 27) {real, imag} */,
  {32'hc22f0106, 32'hc1fbb888} /* (22, 6, 26) {real, imag} */,
  {32'hc28fb56f, 32'h422c2084} /* (22, 6, 25) {real, imag} */,
  {32'h42b3236c, 32'hc28a06ac} /* (22, 6, 24) {real, imag} */,
  {32'hc24f3d2e, 32'h419f19ec} /* (22, 6, 23) {real, imag} */,
  {32'hc2a81e30, 32'h421f150c} /* (22, 6, 22) {real, imag} */,
  {32'h3f1a51c0, 32'h402c2fb0} /* (22, 6, 21) {real, imag} */,
  {32'hc21bd3c8, 32'hc2b9742a} /* (22, 6, 20) {real, imag} */,
  {32'h42d697ce, 32'hc1e7fc09} /* (22, 6, 19) {real, imag} */,
  {32'hbfae0818, 32'hc084ee60} /* (22, 6, 18) {real, imag} */,
  {32'h3f495b90, 32'h428006e0} /* (22, 6, 17) {real, imag} */,
  {32'hc22c40c6, 32'h00000000} /* (22, 6, 16) {real, imag} */,
  {32'h3f495b90, 32'hc28006e0} /* (22, 6, 15) {real, imag} */,
  {32'hbfae0818, 32'h4084ee60} /* (22, 6, 14) {real, imag} */,
  {32'h42d697ce, 32'h41e7fc09} /* (22, 6, 13) {real, imag} */,
  {32'hc21bd3c8, 32'h42b9742a} /* (22, 6, 12) {real, imag} */,
  {32'h3f1a51c0, 32'hc02c2fb0} /* (22, 6, 11) {real, imag} */,
  {32'hc2a81e30, 32'hc21f150c} /* (22, 6, 10) {real, imag} */,
  {32'hc24f3d2e, 32'hc19f19ec} /* (22, 6, 9) {real, imag} */,
  {32'h42b3236c, 32'h428a06ac} /* (22, 6, 8) {real, imag} */,
  {32'hc28fb56f, 32'hc22c2084} /* (22, 6, 7) {real, imag} */,
  {32'hc22f0106, 32'h41fbb888} /* (22, 6, 6) {real, imag} */,
  {32'h43041655, 32'h429f6f6f} /* (22, 6, 5) {real, imag} */,
  {32'hc2437b90, 32'h42a04fae} /* (22, 6, 4) {real, imag} */,
  {32'h428e0fea, 32'h4155220c} /* (22, 6, 3) {real, imag} */,
  {32'h44476cb4, 32'h44184eec} /* (22, 6, 2) {real, imag} */,
  {32'hc5690f08, 32'hc51c4712} /* (22, 6, 1) {real, imag} */,
  {32'hc58a9bea, 32'h00000000} /* (22, 6, 0) {real, imag} */,
  {32'hc5641607, 32'h454ff2a2} /* (22, 5, 31) {real, imag} */,
  {32'h4350889c, 32'hc43c7ab3} /* (22, 5, 30) {real, imag} */,
  {32'h4320625e, 32'hc2b1f501} /* (22, 5, 29) {real, imag} */,
  {32'h4220f304, 32'hc33f83c5} /* (22, 5, 28) {real, imag} */,
  {32'h4373b8a1, 32'h419e11d4} /* (22, 5, 27) {real, imag} */,
  {32'h4290c0e0, 32'h42388e74} /* (22, 5, 26) {real, imag} */,
  {32'h429cc758, 32'h42efc950} /* (22, 5, 25) {real, imag} */,
  {32'hc2aaeb34, 32'hc29960ba} /* (22, 5, 24) {real, imag} */,
  {32'h431250ee, 32'h4135b392} /* (22, 5, 23) {real, imag} */,
  {32'h41895784, 32'h42f3ba38} /* (22, 5, 22) {real, imag} */,
  {32'h3f8e3dc0, 32'hc20c5b53} /* (22, 5, 21) {real, imag} */,
  {32'hc23ba7d2, 32'hc280954f} /* (22, 5, 20) {real, imag} */,
  {32'hc20277f7, 32'hc1a0965c} /* (22, 5, 19) {real, imag} */,
  {32'hc2b7f611, 32'hc1f69c17} /* (22, 5, 18) {real, imag} */,
  {32'hc1437558, 32'hc2b1b1bc} /* (22, 5, 17) {real, imag} */,
  {32'h41502ccd, 32'h00000000} /* (22, 5, 16) {real, imag} */,
  {32'hc1437558, 32'h42b1b1bc} /* (22, 5, 15) {real, imag} */,
  {32'hc2b7f611, 32'h41f69c17} /* (22, 5, 14) {real, imag} */,
  {32'hc20277f7, 32'h41a0965c} /* (22, 5, 13) {real, imag} */,
  {32'hc23ba7d2, 32'h4280954f} /* (22, 5, 12) {real, imag} */,
  {32'h3f8e3dc0, 32'h420c5b53} /* (22, 5, 11) {real, imag} */,
  {32'h41895784, 32'hc2f3ba38} /* (22, 5, 10) {real, imag} */,
  {32'h431250ee, 32'hc135b392} /* (22, 5, 9) {real, imag} */,
  {32'hc2aaeb34, 32'h429960ba} /* (22, 5, 8) {real, imag} */,
  {32'h429cc758, 32'hc2efc950} /* (22, 5, 7) {real, imag} */,
  {32'h4290c0e0, 32'hc2388e74} /* (22, 5, 6) {real, imag} */,
  {32'h4373b8a1, 32'hc19e11d4} /* (22, 5, 5) {real, imag} */,
  {32'h4220f304, 32'h433f83c5} /* (22, 5, 4) {real, imag} */,
  {32'h4320625e, 32'h42b1f501} /* (22, 5, 3) {real, imag} */,
  {32'h4350889c, 32'h443c7ab3} /* (22, 5, 2) {real, imag} */,
  {32'hc5641607, 32'hc54ff2a2} /* (22, 5, 1) {real, imag} */,
  {32'hc59abef4, 32'h00000000} /* (22, 5, 0) {real, imag} */,
  {32'hc55f1e4f, 32'h4573dcd3} /* (22, 4, 31) {real, imag} */,
  {32'hc354e340, 32'hc455939c} /* (22, 4, 30) {real, imag} */,
  {32'h43692c63, 32'hc309acce} /* (22, 4, 29) {real, imag} */,
  {32'h434732d8, 32'hc37193f9} /* (22, 4, 28) {real, imag} */,
  {32'h43198a63, 32'h42f78426} /* (22, 4, 27) {real, imag} */,
  {32'hc218841d, 32'h4195afd0} /* (22, 4, 26) {real, imag} */,
  {32'h42357918, 32'h40d175e0} /* (22, 4, 25) {real, imag} */,
  {32'hc2898764, 32'h4193b1e4} /* (22, 4, 24) {real, imag} */,
  {32'h42768cdd, 32'h4195d0a6} /* (22, 4, 23) {real, imag} */,
  {32'hc2585294, 32'hc2670a99} /* (22, 4, 22) {real, imag} */,
  {32'h428a7e1d, 32'hc295ee79} /* (22, 4, 21) {real, imag} */,
  {32'hc21ba5e9, 32'h41ec7026} /* (22, 4, 20) {real, imag} */,
  {32'hc273481d, 32'h427595bb} /* (22, 4, 19) {real, imag} */,
  {32'hc231713d, 32'hc199e9b4} /* (22, 4, 18) {real, imag} */,
  {32'h423025be, 32'hbfc12a80} /* (22, 4, 17) {real, imag} */,
  {32'h409a08bc, 32'h00000000} /* (22, 4, 16) {real, imag} */,
  {32'h423025be, 32'h3fc12a80} /* (22, 4, 15) {real, imag} */,
  {32'hc231713d, 32'h4199e9b4} /* (22, 4, 14) {real, imag} */,
  {32'hc273481d, 32'hc27595bb} /* (22, 4, 13) {real, imag} */,
  {32'hc21ba5e9, 32'hc1ec7026} /* (22, 4, 12) {real, imag} */,
  {32'h428a7e1d, 32'h4295ee79} /* (22, 4, 11) {real, imag} */,
  {32'hc2585294, 32'h42670a99} /* (22, 4, 10) {real, imag} */,
  {32'h42768cdd, 32'hc195d0a6} /* (22, 4, 9) {real, imag} */,
  {32'hc2898764, 32'hc193b1e4} /* (22, 4, 8) {real, imag} */,
  {32'h42357918, 32'hc0d175e0} /* (22, 4, 7) {real, imag} */,
  {32'hc218841d, 32'hc195afd0} /* (22, 4, 6) {real, imag} */,
  {32'h43198a63, 32'hc2f78426} /* (22, 4, 5) {real, imag} */,
  {32'h434732d8, 32'h437193f9} /* (22, 4, 4) {real, imag} */,
  {32'h43692c63, 32'h4309acce} /* (22, 4, 3) {real, imag} */,
  {32'hc354e340, 32'h4455939c} /* (22, 4, 2) {real, imag} */,
  {32'hc55f1e4f, 32'hc573dcd3} /* (22, 4, 1) {real, imag} */,
  {32'hc5a1a571, 32'h00000000} /* (22, 4, 0) {real, imag} */,
  {32'hc563230c, 32'h457d6a7c} /* (22, 3, 31) {real, imag} */,
  {32'hc38b77ca, 32'hc480e984} /* (22, 3, 30) {real, imag} */,
  {32'h4371119b, 32'hc360de58} /* (22, 3, 29) {real, imag} */,
  {32'h431c62e2, 32'hc3ad30fd} /* (22, 3, 28) {real, imag} */,
  {32'h439c4fc4, 32'h41cc30d8} /* (22, 3, 27) {real, imag} */,
  {32'hc1921fec, 32'hc254e9c7} /* (22, 3, 26) {real, imag} */,
  {32'h4256bf5f, 32'h430af6fa} /* (22, 3, 25) {real, imag} */,
  {32'hc2ae6820, 32'hc2087a4a} /* (22, 3, 24) {real, imag} */,
  {32'h42d13f5f, 32'hc20dd242} /* (22, 3, 23) {real, imag} */,
  {32'h428c982c, 32'hc148e0f3} /* (22, 3, 22) {real, imag} */,
  {32'hc1dfb67c, 32'h420c29da} /* (22, 3, 21) {real, imag} */,
  {32'h42ab828f, 32'h41d3d21d} /* (22, 3, 20) {real, imag} */,
  {32'hc298c91a, 32'hc28d8388} /* (22, 3, 19) {real, imag} */,
  {32'hc2f75136, 32'h4228d112} /* (22, 3, 18) {real, imag} */,
  {32'hc1d2f124, 32'h424ae9a0} /* (22, 3, 17) {real, imag} */,
  {32'h42a1c122, 32'h00000000} /* (22, 3, 16) {real, imag} */,
  {32'hc1d2f124, 32'hc24ae9a0} /* (22, 3, 15) {real, imag} */,
  {32'hc2f75136, 32'hc228d112} /* (22, 3, 14) {real, imag} */,
  {32'hc298c91a, 32'h428d8388} /* (22, 3, 13) {real, imag} */,
  {32'h42ab828f, 32'hc1d3d21d} /* (22, 3, 12) {real, imag} */,
  {32'hc1dfb67c, 32'hc20c29da} /* (22, 3, 11) {real, imag} */,
  {32'h428c982c, 32'h4148e0f3} /* (22, 3, 10) {real, imag} */,
  {32'h42d13f5f, 32'h420dd242} /* (22, 3, 9) {real, imag} */,
  {32'hc2ae6820, 32'h42087a4a} /* (22, 3, 8) {real, imag} */,
  {32'h4256bf5f, 32'hc30af6fa} /* (22, 3, 7) {real, imag} */,
  {32'hc1921fec, 32'h4254e9c7} /* (22, 3, 6) {real, imag} */,
  {32'h439c4fc4, 32'hc1cc30d8} /* (22, 3, 5) {real, imag} */,
  {32'h431c62e2, 32'h43ad30fd} /* (22, 3, 4) {real, imag} */,
  {32'h4371119b, 32'h4360de58} /* (22, 3, 3) {real, imag} */,
  {32'hc38b77ca, 32'h4480e984} /* (22, 3, 2) {real, imag} */,
  {32'hc563230c, 32'hc57d6a7c} /* (22, 3, 1) {real, imag} */,
  {32'hc5ad2dd0, 32'h00000000} /* (22, 3, 0) {real, imag} */,
  {32'hc55e5e92, 32'h45735cd5} /* (22, 2, 31) {real, imag} */,
  {32'hc3ab9b2c, 32'hc4601c42} /* (22, 2, 30) {real, imag} */,
  {32'h428fb063, 32'hc2c5ffea} /* (22, 2, 29) {real, imag} */,
  {32'h42a2327c, 32'hc3922c77} /* (22, 2, 28) {real, imag} */,
  {32'h43876cdd, 32'h42dabcc9} /* (22, 2, 27) {real, imag} */,
  {32'h426a5c8d, 32'hc2cef329} /* (22, 2, 26) {real, imag} */,
  {32'h42da964c, 32'hc2885e51} /* (22, 2, 25) {real, imag} */,
  {32'h4211654c, 32'hc26ceb3e} /* (22, 2, 24) {real, imag} */,
  {32'h4306ab7b, 32'hc24ddad2} /* (22, 2, 23) {real, imag} */,
  {32'hc093d148, 32'hc2858c76} /* (22, 2, 22) {real, imag} */,
  {32'h424295aa, 32'hc22c0174} /* (22, 2, 21) {real, imag} */,
  {32'h4264baa7, 32'h42b06548} /* (22, 2, 20) {real, imag} */,
  {32'hc11cb1e6, 32'hc183dfd3} /* (22, 2, 19) {real, imag} */,
  {32'h40959b94, 32'h3ea10b80} /* (22, 2, 18) {real, imag} */,
  {32'hc12b7dc6, 32'h42295231} /* (22, 2, 17) {real, imag} */,
  {32'h42a9de29, 32'h00000000} /* (22, 2, 16) {real, imag} */,
  {32'hc12b7dc6, 32'hc2295231} /* (22, 2, 15) {real, imag} */,
  {32'h40959b94, 32'hbea10b80} /* (22, 2, 14) {real, imag} */,
  {32'hc11cb1e6, 32'h4183dfd3} /* (22, 2, 13) {real, imag} */,
  {32'h4264baa7, 32'hc2b06548} /* (22, 2, 12) {real, imag} */,
  {32'h424295aa, 32'h422c0174} /* (22, 2, 11) {real, imag} */,
  {32'hc093d148, 32'h42858c76} /* (22, 2, 10) {real, imag} */,
  {32'h4306ab7b, 32'h424ddad2} /* (22, 2, 9) {real, imag} */,
  {32'h4211654c, 32'h426ceb3e} /* (22, 2, 8) {real, imag} */,
  {32'h42da964c, 32'h42885e51} /* (22, 2, 7) {real, imag} */,
  {32'h426a5c8d, 32'h42cef329} /* (22, 2, 6) {real, imag} */,
  {32'h43876cdd, 32'hc2dabcc9} /* (22, 2, 5) {real, imag} */,
  {32'h42a2327c, 32'h43922c77} /* (22, 2, 4) {real, imag} */,
  {32'h428fb063, 32'h42c5ffea} /* (22, 2, 3) {real, imag} */,
  {32'hc3ab9b2c, 32'h44601c42} /* (22, 2, 2) {real, imag} */,
  {32'hc55e5e92, 32'hc5735cd5} /* (22, 2, 1) {real, imag} */,
  {32'hc5ae534f, 32'h00000000} /* (22, 2, 0) {real, imag} */,
  {32'hc5578861, 32'h4564a5ac} /* (22, 1, 31) {real, imag} */,
  {32'hc30d3774, 32'hc455ec82} /* (22, 1, 30) {real, imag} */,
  {32'h431abde9, 32'hc301e0da} /* (22, 1, 29) {real, imag} */,
  {32'h41721e50, 32'hc3b6c2ae} /* (22, 1, 28) {real, imag} */,
  {32'h4345f4b9, 32'h431b846f} /* (22, 1, 27) {real, imag} */,
  {32'hc25d97bc, 32'hc2203372} /* (22, 1, 26) {real, imag} */,
  {32'h42e10d4a, 32'h4227f504} /* (22, 1, 25) {real, imag} */,
  {32'h41505c9a, 32'hc242a7f2} /* (22, 1, 24) {real, imag} */,
  {32'h418b5d4e, 32'hc155949d} /* (22, 1, 23) {real, imag} */,
  {32'hc2a4b6a0, 32'hc163ca42} /* (22, 1, 22) {real, imag} */,
  {32'h41240409, 32'h4254fa5c} /* (22, 1, 21) {real, imag} */,
  {32'h4291a950, 32'hc088e200} /* (22, 1, 20) {real, imag} */,
  {32'hc192821e, 32'h41b993a7} /* (22, 1, 19) {real, imag} */,
  {32'h41a809dc, 32'h405a7bb8} /* (22, 1, 18) {real, imag} */,
  {32'hc2664644, 32'h3fa11d8e} /* (22, 1, 17) {real, imag} */,
  {32'h40a2981e, 32'h00000000} /* (22, 1, 16) {real, imag} */,
  {32'hc2664644, 32'hbfa11d8e} /* (22, 1, 15) {real, imag} */,
  {32'h41a809dc, 32'hc05a7bb8} /* (22, 1, 14) {real, imag} */,
  {32'hc192821e, 32'hc1b993a7} /* (22, 1, 13) {real, imag} */,
  {32'h4291a950, 32'h4088e200} /* (22, 1, 12) {real, imag} */,
  {32'h41240409, 32'hc254fa5c} /* (22, 1, 11) {real, imag} */,
  {32'hc2a4b6a0, 32'h4163ca42} /* (22, 1, 10) {real, imag} */,
  {32'h418b5d4e, 32'h4155949d} /* (22, 1, 9) {real, imag} */,
  {32'h41505c9a, 32'h4242a7f2} /* (22, 1, 8) {real, imag} */,
  {32'h42e10d4a, 32'hc227f504} /* (22, 1, 7) {real, imag} */,
  {32'hc25d97bc, 32'h42203372} /* (22, 1, 6) {real, imag} */,
  {32'h4345f4b9, 32'hc31b846f} /* (22, 1, 5) {real, imag} */,
  {32'h41721e50, 32'h43b6c2ae} /* (22, 1, 4) {real, imag} */,
  {32'h431abde9, 32'h4301e0da} /* (22, 1, 3) {real, imag} */,
  {32'hc30d3774, 32'h4455ec82} /* (22, 1, 2) {real, imag} */,
  {32'hc5578861, 32'hc564a5ac} /* (22, 1, 1) {real, imag} */,
  {32'hc5aaf37d, 32'h00000000} /* (22, 1, 0) {real, imag} */,
  {32'hc563ca4d, 32'h453b8352} /* (22, 0, 31) {real, imag} */,
  {32'h4367a458, 32'hc41e11ca} /* (22, 0, 30) {real, imag} */,
  {32'h43235c11, 32'hc1e33c44} /* (22, 0, 29) {real, imag} */,
  {32'hc260803c, 32'hc36e554d} /* (22, 0, 28) {real, imag} */,
  {32'h417f1aa0, 32'hc1cf3cc4} /* (22, 0, 27) {real, imag} */,
  {32'hc2c62a22, 32'h415c7758} /* (22, 0, 26) {real, imag} */,
  {32'h4226340f, 32'h4230ba3e} /* (22, 0, 25) {real, imag} */,
  {32'h41dbb023, 32'hc28d8ca3} /* (22, 0, 24) {real, imag} */,
  {32'h42873d71, 32'hc2a4a704} /* (22, 0, 23) {real, imag} */,
  {32'hc309fc32, 32'hc2a8e122} /* (22, 0, 22) {real, imag} */,
  {32'hc1f979b8, 32'h41f439de} /* (22, 0, 21) {real, imag} */,
  {32'h422f6ada, 32'h4231f776} /* (22, 0, 20) {real, imag} */,
  {32'hc251cc98, 32'hc27628d0} /* (22, 0, 19) {real, imag} */,
  {32'h423bb08e, 32'h4146ba43} /* (22, 0, 18) {real, imag} */,
  {32'hc104c146, 32'hc2786220} /* (22, 0, 17) {real, imag} */,
  {32'hc25c3935, 32'h00000000} /* (22, 0, 16) {real, imag} */,
  {32'hc104c146, 32'h42786220} /* (22, 0, 15) {real, imag} */,
  {32'h423bb08e, 32'hc146ba43} /* (22, 0, 14) {real, imag} */,
  {32'hc251cc98, 32'h427628d0} /* (22, 0, 13) {real, imag} */,
  {32'h422f6ada, 32'hc231f776} /* (22, 0, 12) {real, imag} */,
  {32'hc1f979b8, 32'hc1f439de} /* (22, 0, 11) {real, imag} */,
  {32'hc309fc32, 32'h42a8e122} /* (22, 0, 10) {real, imag} */,
  {32'h42873d71, 32'h42a4a704} /* (22, 0, 9) {real, imag} */,
  {32'h41dbb023, 32'h428d8ca3} /* (22, 0, 8) {real, imag} */,
  {32'h4226340f, 32'hc230ba3e} /* (22, 0, 7) {real, imag} */,
  {32'hc2c62a22, 32'hc15c7758} /* (22, 0, 6) {real, imag} */,
  {32'h417f1aa0, 32'h41cf3cc4} /* (22, 0, 5) {real, imag} */,
  {32'hc260803c, 32'h436e554d} /* (22, 0, 4) {real, imag} */,
  {32'h43235c11, 32'h41e33c44} /* (22, 0, 3) {real, imag} */,
  {32'h4367a458, 32'h441e11ca} /* (22, 0, 2) {real, imag} */,
  {32'hc563ca4d, 32'hc53b8352} /* (22, 0, 1) {real, imag} */,
  {32'hc5a5510d, 32'h00000000} /* (22, 0, 0) {real, imag} */,
  {32'hc583f146, 32'h4515235c} /* (21, 31, 31) {real, imag} */,
  {32'h4447e62b, 32'hc4040067} /* (21, 31, 30) {real, imag} */,
  {32'h41dd09b8, 32'h4277b55c} /* (21, 31, 29) {real, imag} */,
  {32'hc2de38ed, 32'hc20f3da0} /* (21, 31, 28) {real, imag} */,
  {32'h42410f80, 32'hc1a538e6} /* (21, 31, 27) {real, imag} */,
  {32'h413d54a8, 32'hc245a486} /* (21, 31, 26) {real, imag} */,
  {32'h4298a9fb, 32'h41b82382} /* (21, 31, 25) {real, imag} */,
  {32'h4209b68a, 32'h40074518} /* (21, 31, 24) {real, imag} */,
  {32'hbca49000, 32'h4245ba37} /* (21, 31, 23) {real, imag} */,
  {32'h415bbbf4, 32'h41e1a820} /* (21, 31, 22) {real, imag} */,
  {32'h41779bd8, 32'hc28f7a23} /* (21, 31, 21) {real, imag} */,
  {32'h4239f976, 32'hc1c716dc} /* (21, 31, 20) {real, imag} */,
  {32'hc17d1262, 32'h41992f46} /* (21, 31, 19) {real, imag} */,
  {32'hc229faec, 32'hc18eed1e} /* (21, 31, 18) {real, imag} */,
  {32'hc11123bb, 32'hc1d32df3} /* (21, 31, 17) {real, imag} */,
  {32'h42000ee4, 32'h00000000} /* (21, 31, 16) {real, imag} */,
  {32'hc11123bb, 32'h41d32df3} /* (21, 31, 15) {real, imag} */,
  {32'hc229faec, 32'h418eed1e} /* (21, 31, 14) {real, imag} */,
  {32'hc17d1262, 32'hc1992f46} /* (21, 31, 13) {real, imag} */,
  {32'h4239f976, 32'h41c716dc} /* (21, 31, 12) {real, imag} */,
  {32'h41779bd8, 32'h428f7a23} /* (21, 31, 11) {real, imag} */,
  {32'h415bbbf4, 32'hc1e1a820} /* (21, 31, 10) {real, imag} */,
  {32'hbca49000, 32'hc245ba37} /* (21, 31, 9) {real, imag} */,
  {32'h4209b68a, 32'hc0074518} /* (21, 31, 8) {real, imag} */,
  {32'h4298a9fb, 32'hc1b82382} /* (21, 31, 7) {real, imag} */,
  {32'h413d54a8, 32'h4245a486} /* (21, 31, 6) {real, imag} */,
  {32'h42410f80, 32'h41a538e6} /* (21, 31, 5) {real, imag} */,
  {32'hc2de38ed, 32'h420f3da0} /* (21, 31, 4) {real, imag} */,
  {32'h41dd09b8, 32'hc277b55c} /* (21, 31, 3) {real, imag} */,
  {32'h4447e62b, 32'h44040067} /* (21, 31, 2) {real, imag} */,
  {32'hc583f146, 32'hc515235c} /* (21, 31, 1) {real, imag} */,
  {32'hc5a6ed23, 32'h00000000} /* (21, 31, 0) {real, imag} */,
  {32'hc5967bf2, 32'h4501178e} /* (21, 30, 31) {real, imag} */,
  {32'h4491c5ce, 32'hc3fd97cc} /* (21, 30, 30) {real, imag} */,
  {32'hc1cf4c4c, 32'h423878aa} /* (21, 30, 29) {real, imag} */,
  {32'hc38abaf4, 32'h40e51d80} /* (21, 30, 28) {real, imag} */,
  {32'h43522419, 32'hc28ed907} /* (21, 30, 27) {real, imag} */,
  {32'hc3034682, 32'hc31f7dfa} /* (21, 30, 26) {real, imag} */,
  {32'h41a7cabe, 32'h420e0754} /* (21, 30, 25) {real, imag} */,
  {32'h4273ddaa, 32'hc2bd5efa} /* (21, 30, 24) {real, imag} */,
  {32'h42390803, 32'hc10d5406} /* (21, 30, 23) {real, imag} */,
  {32'h41edf2f6, 32'h42978160} /* (21, 30, 22) {real, imag} */,
  {32'h41c38786, 32'h4134aa74} /* (21, 30, 21) {real, imag} */,
  {32'h42f27eee, 32'hc2a4b384} /* (21, 30, 20) {real, imag} */,
  {32'hc22ea698, 32'hc1c2ca76} /* (21, 30, 19) {real, imag} */,
  {32'h4244169e, 32'h4223deee} /* (21, 30, 18) {real, imag} */,
  {32'h41e34f22, 32'hc20e7902} /* (21, 30, 17) {real, imag} */,
  {32'hc1d44e4b, 32'h00000000} /* (21, 30, 16) {real, imag} */,
  {32'h41e34f22, 32'h420e7902} /* (21, 30, 15) {real, imag} */,
  {32'h4244169e, 32'hc223deee} /* (21, 30, 14) {real, imag} */,
  {32'hc22ea698, 32'h41c2ca76} /* (21, 30, 13) {real, imag} */,
  {32'h42f27eee, 32'h42a4b384} /* (21, 30, 12) {real, imag} */,
  {32'h41c38786, 32'hc134aa74} /* (21, 30, 11) {real, imag} */,
  {32'h41edf2f6, 32'hc2978160} /* (21, 30, 10) {real, imag} */,
  {32'h42390803, 32'h410d5406} /* (21, 30, 9) {real, imag} */,
  {32'h4273ddaa, 32'h42bd5efa} /* (21, 30, 8) {real, imag} */,
  {32'h41a7cabe, 32'hc20e0754} /* (21, 30, 7) {real, imag} */,
  {32'hc3034682, 32'h431f7dfa} /* (21, 30, 6) {real, imag} */,
  {32'h43522419, 32'h428ed907} /* (21, 30, 5) {real, imag} */,
  {32'hc38abaf4, 32'hc0e51d80} /* (21, 30, 4) {real, imag} */,
  {32'hc1cf4c4c, 32'hc23878aa} /* (21, 30, 3) {real, imag} */,
  {32'h4491c5ce, 32'h43fd97cc} /* (21, 30, 2) {real, imag} */,
  {32'hc5967bf2, 32'hc501178e} /* (21, 30, 1) {real, imag} */,
  {32'hc5a8a248, 32'h00000000} /* (21, 30, 0) {real, imag} */,
  {32'hc5a5df93, 32'h44cada0f} /* (21, 29, 31) {real, imag} */,
  {32'h44b96039, 32'hc3925047} /* (21, 29, 30) {real, imag} */,
  {32'hc1e6ddc8, 32'hc2a680f9} /* (21, 29, 29) {real, imag} */,
  {32'hc3ada238, 32'h4316d57a} /* (21, 29, 28) {real, imag} */,
  {32'h43828922, 32'hc29af5b4} /* (21, 29, 27) {real, imag} */,
  {32'h4186600d, 32'h42503f88} /* (21, 29, 26) {real, imag} */,
  {32'h4001020c, 32'h421b4047} /* (21, 29, 25) {real, imag} */,
  {32'h42a1b061, 32'hc23dd0a3} /* (21, 29, 24) {real, imag} */,
  {32'h4269278e, 32'hc0b74d68} /* (21, 29, 23) {real, imag} */,
  {32'h425f1bea, 32'h40595ce4} /* (21, 29, 22) {real, imag} */,
  {32'h42dafa8b, 32'h41a64624} /* (21, 29, 21) {real, imag} */,
  {32'h425e68f6, 32'hc2f806b7} /* (21, 29, 20) {real, imag} */,
  {32'h4216a31a, 32'hc198457a} /* (21, 29, 19) {real, imag} */,
  {32'hbec4f780, 32'hc22b247b} /* (21, 29, 18) {real, imag} */,
  {32'hc204588e, 32'h41aa0f90} /* (21, 29, 17) {real, imag} */,
  {32'h428a2aa9, 32'h00000000} /* (21, 29, 16) {real, imag} */,
  {32'hc204588e, 32'hc1aa0f90} /* (21, 29, 15) {real, imag} */,
  {32'hbec4f780, 32'h422b247b} /* (21, 29, 14) {real, imag} */,
  {32'h4216a31a, 32'h4198457a} /* (21, 29, 13) {real, imag} */,
  {32'h425e68f6, 32'h42f806b7} /* (21, 29, 12) {real, imag} */,
  {32'h42dafa8b, 32'hc1a64624} /* (21, 29, 11) {real, imag} */,
  {32'h425f1bea, 32'hc0595ce4} /* (21, 29, 10) {real, imag} */,
  {32'h4269278e, 32'h40b74d68} /* (21, 29, 9) {real, imag} */,
  {32'h42a1b061, 32'h423dd0a3} /* (21, 29, 8) {real, imag} */,
  {32'h4001020c, 32'hc21b4047} /* (21, 29, 7) {real, imag} */,
  {32'h4186600d, 32'hc2503f88} /* (21, 29, 6) {real, imag} */,
  {32'h43828922, 32'h429af5b4} /* (21, 29, 5) {real, imag} */,
  {32'hc3ada238, 32'hc316d57a} /* (21, 29, 4) {real, imag} */,
  {32'hc1e6ddc8, 32'h42a680f9} /* (21, 29, 3) {real, imag} */,
  {32'h44b96039, 32'h43925047} /* (21, 29, 2) {real, imag} */,
  {32'hc5a5df93, 32'hc4cada0f} /* (21, 29, 1) {real, imag} */,
  {32'hc5a9a986, 32'h00000000} /* (21, 29, 0) {real, imag} */,
  {32'hc5ab00b6, 32'h44a98c96} /* (21, 28, 31) {real, imag} */,
  {32'h44e4d8ac, 32'hc3e9d5b4} /* (21, 28, 30) {real, imag} */,
  {32'hc1ffaeb0, 32'hc1a5ebbc} /* (21, 28, 29) {real, imag} */,
  {32'hc38c686e, 32'h4324dfbe} /* (21, 28, 28) {real, imag} */,
  {32'h4360a86a, 32'hc345ca52} /* (21, 28, 27) {real, imag} */,
  {32'hc205e580, 32'h42495d4f} /* (21, 28, 26) {real, imag} */,
  {32'hc2ea3b88, 32'h42949646} /* (21, 28, 25) {real, imag} */,
  {32'hc07d48e0, 32'hc2d7bb48} /* (21, 28, 24) {real, imag} */,
  {32'hc196e03e, 32'h42afcc20} /* (21, 28, 23) {real, imag} */,
  {32'hc2849bb5, 32'hc1923150} /* (21, 28, 22) {real, imag} */,
  {32'h4202242c, 32'hc2c90f1a} /* (21, 28, 21) {real, imag} */,
  {32'h41f6bc80, 32'hc29491b3} /* (21, 28, 20) {real, imag} */,
  {32'hc222912b, 32'hc2c9ee7a} /* (21, 28, 19) {real, imag} */,
  {32'hc2ca01b6, 32'h41f88950} /* (21, 28, 18) {real, imag} */,
  {32'hc27451c6, 32'hc163dfb3} /* (21, 28, 17) {real, imag} */,
  {32'h42c51e36, 32'h00000000} /* (21, 28, 16) {real, imag} */,
  {32'hc27451c6, 32'h4163dfb3} /* (21, 28, 15) {real, imag} */,
  {32'hc2ca01b6, 32'hc1f88950} /* (21, 28, 14) {real, imag} */,
  {32'hc222912b, 32'h42c9ee7a} /* (21, 28, 13) {real, imag} */,
  {32'h41f6bc80, 32'h429491b3} /* (21, 28, 12) {real, imag} */,
  {32'h4202242c, 32'h42c90f1a} /* (21, 28, 11) {real, imag} */,
  {32'hc2849bb5, 32'h41923150} /* (21, 28, 10) {real, imag} */,
  {32'hc196e03e, 32'hc2afcc20} /* (21, 28, 9) {real, imag} */,
  {32'hc07d48e0, 32'h42d7bb48} /* (21, 28, 8) {real, imag} */,
  {32'hc2ea3b88, 32'hc2949646} /* (21, 28, 7) {real, imag} */,
  {32'hc205e580, 32'hc2495d4f} /* (21, 28, 6) {real, imag} */,
  {32'h4360a86a, 32'h4345ca52} /* (21, 28, 5) {real, imag} */,
  {32'hc38c686e, 32'hc324dfbe} /* (21, 28, 4) {real, imag} */,
  {32'hc1ffaeb0, 32'h41a5ebbc} /* (21, 28, 3) {real, imag} */,
  {32'h44e4d8ac, 32'h43e9d5b4} /* (21, 28, 2) {real, imag} */,
  {32'hc5ab00b6, 32'hc4a98c96} /* (21, 28, 1) {real, imag} */,
  {32'hc5b4669b, 32'h00000000} /* (21, 28, 0) {real, imag} */,
  {32'hc5a9521a, 32'h44929c13} /* (21, 27, 31) {real, imag} */,
  {32'h44eada86, 32'hc4027ef1} /* (21, 27, 30) {real, imag} */,
  {32'hc10bd296, 32'h405e1ca0} /* (21, 27, 29) {real, imag} */,
  {32'hc370cfe4, 32'h42894972} /* (21, 27, 28) {real, imag} */,
  {32'h4345d038, 32'hc334a808} /* (21, 27, 27) {real, imag} */,
  {32'hc22cb339, 32'hc31ddf3f} /* (21, 27, 26) {real, imag} */,
  {32'hc2c0b8bf, 32'hc0661890} /* (21, 27, 25) {real, imag} */,
  {32'h41b28eaf, 32'hc23804a9} /* (21, 27, 24) {real, imag} */,
  {32'h42b16636, 32'h411f7c4f} /* (21, 27, 23) {real, imag} */,
  {32'hc2013311, 32'h41c5a20e} /* (21, 27, 22) {real, imag} */,
  {32'h42669882, 32'h42811c14} /* (21, 27, 21) {real, imag} */,
  {32'hc279b1d6, 32'h41cfd993} /* (21, 27, 20) {real, imag} */,
  {32'h409605e0, 32'h41b10704} /* (21, 27, 19) {real, imag} */,
  {32'h4235389c, 32'h414a2b3c} /* (21, 27, 18) {real, imag} */,
  {32'hc02fc074, 32'h421d9ba4} /* (21, 27, 17) {real, imag} */,
  {32'hc312b8a9, 32'h00000000} /* (21, 27, 16) {real, imag} */,
  {32'hc02fc074, 32'hc21d9ba4} /* (21, 27, 15) {real, imag} */,
  {32'h4235389c, 32'hc14a2b3c} /* (21, 27, 14) {real, imag} */,
  {32'h409605e0, 32'hc1b10704} /* (21, 27, 13) {real, imag} */,
  {32'hc279b1d6, 32'hc1cfd993} /* (21, 27, 12) {real, imag} */,
  {32'h42669882, 32'hc2811c14} /* (21, 27, 11) {real, imag} */,
  {32'hc2013311, 32'hc1c5a20e} /* (21, 27, 10) {real, imag} */,
  {32'h42b16636, 32'hc11f7c4f} /* (21, 27, 9) {real, imag} */,
  {32'h41b28eaf, 32'h423804a9} /* (21, 27, 8) {real, imag} */,
  {32'hc2c0b8bf, 32'h40661890} /* (21, 27, 7) {real, imag} */,
  {32'hc22cb339, 32'h431ddf3f} /* (21, 27, 6) {real, imag} */,
  {32'h4345d038, 32'h4334a808} /* (21, 27, 5) {real, imag} */,
  {32'hc370cfe4, 32'hc2894972} /* (21, 27, 4) {real, imag} */,
  {32'hc10bd296, 32'hc05e1ca0} /* (21, 27, 3) {real, imag} */,
  {32'h44eada86, 32'h44027ef1} /* (21, 27, 2) {real, imag} */,
  {32'hc5a9521a, 32'hc4929c13} /* (21, 27, 1) {real, imag} */,
  {32'hc5b9eb55, 32'h00000000} /* (21, 27, 0) {real, imag} */,
  {32'hc5a4d6b2, 32'h4476f4dd} /* (21, 26, 31) {real, imag} */,
  {32'h44f94024, 32'hc3c89274} /* (21, 26, 30) {real, imag} */,
  {32'hc1b1a601, 32'h4121316a} /* (21, 26, 29) {real, imag} */,
  {32'hc3b6c335, 32'h40b0acb0} /* (21, 26, 28) {real, imag} */,
  {32'h43825d06, 32'hc3168607} /* (21, 26, 27) {real, imag} */,
  {32'h42387ef6, 32'h424dfa6c} /* (21, 26, 26) {real, imag} */,
  {32'hc1eb1864, 32'hc2bbeee3} /* (21, 26, 25) {real, imag} */,
  {32'h427b1879, 32'hc040e328} /* (21, 26, 24) {real, imag} */,
  {32'h4273af6a, 32'h42b393fb} /* (21, 26, 23) {real, imag} */,
  {32'h42f23e48, 32'hc2e1a068} /* (21, 26, 22) {real, imag} */,
  {32'hc29d83da, 32'hc36b4bd6} /* (21, 26, 21) {real, imag} */,
  {32'hc235e344, 32'hc21d8eed} /* (21, 26, 20) {real, imag} */,
  {32'hc2045f50, 32'h41c6134d} /* (21, 26, 19) {real, imag} */,
  {32'h4026ef00, 32'h412b0d42} /* (21, 26, 18) {real, imag} */,
  {32'h4130285a, 32'hc1dbf87f} /* (21, 26, 17) {real, imag} */,
  {32'hc195addf, 32'h00000000} /* (21, 26, 16) {real, imag} */,
  {32'h4130285a, 32'h41dbf87f} /* (21, 26, 15) {real, imag} */,
  {32'h4026ef00, 32'hc12b0d42} /* (21, 26, 14) {real, imag} */,
  {32'hc2045f50, 32'hc1c6134d} /* (21, 26, 13) {real, imag} */,
  {32'hc235e344, 32'h421d8eed} /* (21, 26, 12) {real, imag} */,
  {32'hc29d83da, 32'h436b4bd6} /* (21, 26, 11) {real, imag} */,
  {32'h42f23e48, 32'h42e1a068} /* (21, 26, 10) {real, imag} */,
  {32'h4273af6a, 32'hc2b393fb} /* (21, 26, 9) {real, imag} */,
  {32'h427b1879, 32'h4040e328} /* (21, 26, 8) {real, imag} */,
  {32'hc1eb1864, 32'h42bbeee3} /* (21, 26, 7) {real, imag} */,
  {32'h42387ef6, 32'hc24dfa6c} /* (21, 26, 6) {real, imag} */,
  {32'h43825d06, 32'h43168607} /* (21, 26, 5) {real, imag} */,
  {32'hc3b6c335, 32'hc0b0acb0} /* (21, 26, 4) {real, imag} */,
  {32'hc1b1a601, 32'hc121316a} /* (21, 26, 3) {real, imag} */,
  {32'h44f94024, 32'h43c89274} /* (21, 26, 2) {real, imag} */,
  {32'hc5a4d6b2, 32'hc476f4dd} /* (21, 26, 1) {real, imag} */,
  {32'hc5b00a7f, 32'h00000000} /* (21, 26, 0) {real, imag} */,
  {32'hc59c1ad5, 32'h444aa897} /* (21, 25, 31) {real, imag} */,
  {32'h44f2da24, 32'hc3ca8274} /* (21, 25, 30) {real, imag} */,
  {32'hc2a13a00, 32'h419addfe} /* (21, 25, 29) {real, imag} */,
  {32'hc3395ce1, 32'hc29986de} /* (21, 25, 28) {real, imag} */,
  {32'h438b5af2, 32'hc36623be} /* (21, 25, 27) {real, imag} */,
  {32'hc2890a7c, 32'h4234f54d} /* (21, 25, 26) {real, imag} */,
  {32'hc16d1b28, 32'h42ae1cef} /* (21, 25, 25) {real, imag} */,
  {32'h41e2923a, 32'hc2babdee} /* (21, 25, 24) {real, imag} */,
  {32'h428807e4, 32'h42b5db92} /* (21, 25, 23) {real, imag} */,
  {32'hc01c7bf0, 32'h412b72be} /* (21, 25, 22) {real, imag} */,
  {32'h422d8dac, 32'hc2079a9d} /* (21, 25, 21) {real, imag} */,
  {32'hc23aea4a, 32'h4292318e} /* (21, 25, 20) {real, imag} */,
  {32'hc244da92, 32'h426345bb} /* (21, 25, 19) {real, imag} */,
  {32'h41a8f5aa, 32'h41dfc91d} /* (21, 25, 18) {real, imag} */,
  {32'hc1a0000e, 32'hc20ca0dc} /* (21, 25, 17) {real, imag} */,
  {32'hbfb30e20, 32'h00000000} /* (21, 25, 16) {real, imag} */,
  {32'hc1a0000e, 32'h420ca0dc} /* (21, 25, 15) {real, imag} */,
  {32'h41a8f5aa, 32'hc1dfc91d} /* (21, 25, 14) {real, imag} */,
  {32'hc244da92, 32'hc26345bb} /* (21, 25, 13) {real, imag} */,
  {32'hc23aea4a, 32'hc292318e} /* (21, 25, 12) {real, imag} */,
  {32'h422d8dac, 32'h42079a9d} /* (21, 25, 11) {real, imag} */,
  {32'hc01c7bf0, 32'hc12b72be} /* (21, 25, 10) {real, imag} */,
  {32'h428807e4, 32'hc2b5db92} /* (21, 25, 9) {real, imag} */,
  {32'h41e2923a, 32'h42babdee} /* (21, 25, 8) {real, imag} */,
  {32'hc16d1b28, 32'hc2ae1cef} /* (21, 25, 7) {real, imag} */,
  {32'hc2890a7c, 32'hc234f54d} /* (21, 25, 6) {real, imag} */,
  {32'h438b5af2, 32'h436623be} /* (21, 25, 5) {real, imag} */,
  {32'hc3395ce1, 32'h429986de} /* (21, 25, 4) {real, imag} */,
  {32'hc2a13a00, 32'hc19addfe} /* (21, 25, 3) {real, imag} */,
  {32'h44f2da24, 32'h43ca8274} /* (21, 25, 2) {real, imag} */,
  {32'hc59c1ad5, 32'hc44aa897} /* (21, 25, 1) {real, imag} */,
  {32'hc59f28fd, 32'h00000000} /* (21, 25, 0) {real, imag} */,
  {32'hc588f257, 32'h44016d16} /* (21, 24, 31) {real, imag} */,
  {32'h44d5b090, 32'hc3f1ba10} /* (21, 24, 30) {real, imag} */,
  {32'hc28fdbc3, 32'hc268d4e2} /* (21, 24, 29) {real, imag} */,
  {32'hc364e92e, 32'h42e7391f} /* (21, 24, 28) {real, imag} */,
  {32'h437ae9b2, 32'hc347afd9} /* (21, 24, 27) {real, imag} */,
  {32'hc28bdd4a, 32'hc2b1db42} /* (21, 24, 26) {real, imag} */,
  {32'hbfb792d0, 32'h42301d35} /* (21, 24, 25) {real, imag} */,
  {32'h42dd34f4, 32'hc2eb958c} /* (21, 24, 24) {real, imag} */,
  {32'h427ea4d9, 32'h4300b2aa} /* (21, 24, 23) {real, imag} */,
  {32'h41788123, 32'hc28787a1} /* (21, 24, 22) {real, imag} */,
  {32'hc2370dde, 32'h4152f2f6} /* (21, 24, 21) {real, imag} */,
  {32'h4267fbc4, 32'hc19fac0c} /* (21, 24, 20) {real, imag} */,
  {32'h40129070, 32'h42b295ed} /* (21, 24, 19) {real, imag} */,
  {32'h42c91d7f, 32'hc20940c1} /* (21, 24, 18) {real, imag} */,
  {32'hc26b6418, 32'hc1f1e73e} /* (21, 24, 17) {real, imag} */,
  {32'h3ff0a298, 32'h00000000} /* (21, 24, 16) {real, imag} */,
  {32'hc26b6418, 32'h41f1e73e} /* (21, 24, 15) {real, imag} */,
  {32'h42c91d7f, 32'h420940c1} /* (21, 24, 14) {real, imag} */,
  {32'h40129070, 32'hc2b295ed} /* (21, 24, 13) {real, imag} */,
  {32'h4267fbc4, 32'h419fac0c} /* (21, 24, 12) {real, imag} */,
  {32'hc2370dde, 32'hc152f2f6} /* (21, 24, 11) {real, imag} */,
  {32'h41788123, 32'h428787a1} /* (21, 24, 10) {real, imag} */,
  {32'h427ea4d9, 32'hc300b2aa} /* (21, 24, 9) {real, imag} */,
  {32'h42dd34f4, 32'h42eb958c} /* (21, 24, 8) {real, imag} */,
  {32'hbfb792d0, 32'hc2301d35} /* (21, 24, 7) {real, imag} */,
  {32'hc28bdd4a, 32'h42b1db42} /* (21, 24, 6) {real, imag} */,
  {32'h437ae9b2, 32'h4347afd9} /* (21, 24, 5) {real, imag} */,
  {32'hc364e92e, 32'hc2e7391f} /* (21, 24, 4) {real, imag} */,
  {32'hc28fdbc3, 32'h4268d4e2} /* (21, 24, 3) {real, imag} */,
  {32'h44d5b090, 32'h43f1ba10} /* (21, 24, 2) {real, imag} */,
  {32'hc588f257, 32'hc4016d16} /* (21, 24, 1) {real, imag} */,
  {32'hc582342c, 32'h00000000} /* (21, 24, 0) {real, imag} */,
  {32'hc55fa34c, 32'h43c07232} /* (21, 23, 31) {real, imag} */,
  {32'h44a8bf49, 32'hc3bc09aa} /* (21, 23, 30) {real, imag} */,
  {32'hc19ace06, 32'hbecff360} /* (21, 23, 29) {real, imag} */,
  {32'hc2c6c4f6, 32'h42f0af06} /* (21, 23, 28) {real, imag} */,
  {32'h4382f420, 32'hc1f94652} /* (21, 23, 27) {real, imag} */,
  {32'h41de1909, 32'hc17bc308} /* (21, 23, 26) {real, imag} */,
  {32'hc2d6be16, 32'hc13033cc} /* (21, 23, 25) {real, imag} */,
  {32'h4302bf7b, 32'hc26a6573} /* (21, 23, 24) {real, imag} */,
  {32'hc2bbd81a, 32'hc25aa690} /* (21, 23, 23) {real, imag} */,
  {32'hc1bce542, 32'hc2677b78} /* (21, 23, 22) {real, imag} */,
  {32'h4191f4b4, 32'hc2365814} /* (21, 23, 21) {real, imag} */,
  {32'hc1a25cb6, 32'h4166cba2} /* (21, 23, 20) {real, imag} */,
  {32'hc10cf480, 32'h4222950e} /* (21, 23, 19) {real, imag} */,
  {32'hbfdd8a28, 32'hc2d8a56b} /* (21, 23, 18) {real, imag} */,
  {32'hc1fa1334, 32'hc1154af0} /* (21, 23, 17) {real, imag} */,
  {32'h42905d3e, 32'h00000000} /* (21, 23, 16) {real, imag} */,
  {32'hc1fa1334, 32'h41154af0} /* (21, 23, 15) {real, imag} */,
  {32'hbfdd8a28, 32'h42d8a56b} /* (21, 23, 14) {real, imag} */,
  {32'hc10cf480, 32'hc222950e} /* (21, 23, 13) {real, imag} */,
  {32'hc1a25cb6, 32'hc166cba2} /* (21, 23, 12) {real, imag} */,
  {32'h4191f4b4, 32'h42365814} /* (21, 23, 11) {real, imag} */,
  {32'hc1bce542, 32'h42677b78} /* (21, 23, 10) {real, imag} */,
  {32'hc2bbd81a, 32'h425aa690} /* (21, 23, 9) {real, imag} */,
  {32'h4302bf7b, 32'h426a6573} /* (21, 23, 8) {real, imag} */,
  {32'hc2d6be16, 32'h413033cc} /* (21, 23, 7) {real, imag} */,
  {32'h41de1909, 32'h417bc308} /* (21, 23, 6) {real, imag} */,
  {32'h4382f420, 32'h41f94652} /* (21, 23, 5) {real, imag} */,
  {32'hc2c6c4f6, 32'hc2f0af06} /* (21, 23, 4) {real, imag} */,
  {32'hc19ace06, 32'h3ecff360} /* (21, 23, 3) {real, imag} */,
  {32'h44a8bf49, 32'h43bc09aa} /* (21, 23, 2) {real, imag} */,
  {32'hc55fa34c, 32'hc3c07232} /* (21, 23, 1) {real, imag} */,
  {32'hc5603cea, 32'h00000000} /* (21, 23, 0) {real, imag} */,
  {32'hc521986b, 32'h4332bf70} /* (21, 22, 31) {real, imag} */,
  {32'h4454bd0d, 32'hc3bd62ea} /* (21, 22, 30) {real, imag} */,
  {32'hc2213f66, 32'hc12b728c} /* (21, 22, 29) {real, imag} */,
  {32'hc2ebd888, 32'h4279c787} /* (21, 22, 28) {real, imag} */,
  {32'h438e062e, 32'hc2274f77} /* (21, 22, 27) {real, imag} */,
  {32'hc137fe78, 32'hc29028c9} /* (21, 22, 26) {real, imag} */,
  {32'hc1eeb084, 32'h41f51c09} /* (21, 22, 25) {real, imag} */,
  {32'h425a231b, 32'h41b262f0} /* (21, 22, 24) {real, imag} */,
  {32'hc2a9fdaf, 32'h3fd16cb0} /* (21, 22, 23) {real, imag} */,
  {32'h42510c2e, 32'hc2e84e8a} /* (21, 22, 22) {real, imag} */,
  {32'h40e3cc74, 32'hc201def7} /* (21, 22, 21) {real, imag} */,
  {32'hc21f2c52, 32'hc2811056} /* (21, 22, 20) {real, imag} */,
  {32'h41a609f8, 32'hc073976e} /* (21, 22, 19) {real, imag} */,
  {32'h4235380a, 32'hc2ed7952} /* (21, 22, 18) {real, imag} */,
  {32'h3f8d9328, 32'h426302cc} /* (21, 22, 17) {real, imag} */,
  {32'h4226e010, 32'h00000000} /* (21, 22, 16) {real, imag} */,
  {32'h3f8d9328, 32'hc26302cc} /* (21, 22, 15) {real, imag} */,
  {32'h4235380a, 32'h42ed7952} /* (21, 22, 14) {real, imag} */,
  {32'h41a609f8, 32'h4073976e} /* (21, 22, 13) {real, imag} */,
  {32'hc21f2c52, 32'h42811056} /* (21, 22, 12) {real, imag} */,
  {32'h40e3cc74, 32'h4201def7} /* (21, 22, 11) {real, imag} */,
  {32'h42510c2e, 32'h42e84e8a} /* (21, 22, 10) {real, imag} */,
  {32'hc2a9fdaf, 32'hbfd16cb0} /* (21, 22, 9) {real, imag} */,
  {32'h425a231b, 32'hc1b262f0} /* (21, 22, 8) {real, imag} */,
  {32'hc1eeb084, 32'hc1f51c09} /* (21, 22, 7) {real, imag} */,
  {32'hc137fe78, 32'h429028c9} /* (21, 22, 6) {real, imag} */,
  {32'h438e062e, 32'h42274f77} /* (21, 22, 5) {real, imag} */,
  {32'hc2ebd888, 32'hc279c787} /* (21, 22, 4) {real, imag} */,
  {32'hc2213f66, 32'h412b728c} /* (21, 22, 3) {real, imag} */,
  {32'h4454bd0d, 32'h43bd62ea} /* (21, 22, 2) {real, imag} */,
  {32'hc521986b, 32'hc332bf70} /* (21, 22, 1) {real, imag} */,
  {32'hc51fbb0d, 32'h00000000} /* (21, 22, 0) {real, imag} */,
  {32'hc449cc11, 32'h42175ae0} /* (21, 21, 31) {real, imag} */,
  {32'h43018d42, 32'hc34f30ae} /* (21, 21, 30) {real, imag} */,
  {32'hc24f86e2, 32'h426e68c5} /* (21, 21, 29) {real, imag} */,
  {32'hc312aeb5, 32'hc26b3c08} /* (21, 21, 28) {real, imag} */,
  {32'h42469014, 32'hc239ff65} /* (21, 21, 27) {real, imag} */,
  {32'hc2a32c65, 32'hc1a7e82c} /* (21, 21, 26) {real, imag} */,
  {32'hc08a5a1c, 32'hc1272703} /* (21, 21, 25) {real, imag} */,
  {32'h41699070, 32'hc254a416} /* (21, 21, 24) {real, imag} */,
  {32'hc166659f, 32'h4155b8b9} /* (21, 21, 23) {real, imag} */,
  {32'hc2046bc3, 32'hc2c9f851} /* (21, 21, 22) {real, imag} */,
  {32'h404e5020, 32'h404b7420} /* (21, 21, 21) {real, imag} */,
  {32'h420e4eb8, 32'hc18d94f3} /* (21, 21, 20) {real, imag} */,
  {32'hc042d340, 32'hc2075237} /* (21, 21, 19) {real, imag} */,
  {32'h4218f72b, 32'hc2964e39} /* (21, 21, 18) {real, imag} */,
  {32'h42b3962e, 32'hbfe35a68} /* (21, 21, 17) {real, imag} */,
  {32'hc19aa541, 32'h00000000} /* (21, 21, 16) {real, imag} */,
  {32'h42b3962e, 32'h3fe35a68} /* (21, 21, 15) {real, imag} */,
  {32'h4218f72b, 32'h42964e39} /* (21, 21, 14) {real, imag} */,
  {32'hc042d340, 32'h42075237} /* (21, 21, 13) {real, imag} */,
  {32'h420e4eb8, 32'h418d94f3} /* (21, 21, 12) {real, imag} */,
  {32'h404e5020, 32'hc04b7420} /* (21, 21, 11) {real, imag} */,
  {32'hc2046bc3, 32'h42c9f851} /* (21, 21, 10) {real, imag} */,
  {32'hc166659f, 32'hc155b8b9} /* (21, 21, 9) {real, imag} */,
  {32'h41699070, 32'h4254a416} /* (21, 21, 8) {real, imag} */,
  {32'hc08a5a1c, 32'h41272703} /* (21, 21, 7) {real, imag} */,
  {32'hc2a32c65, 32'h41a7e82c} /* (21, 21, 6) {real, imag} */,
  {32'h42469014, 32'h4239ff65} /* (21, 21, 5) {real, imag} */,
  {32'hc312aeb5, 32'h426b3c08} /* (21, 21, 4) {real, imag} */,
  {32'hc24f86e2, 32'hc26e68c5} /* (21, 21, 3) {real, imag} */,
  {32'h43018d42, 32'h434f30ae} /* (21, 21, 2) {real, imag} */,
  {32'hc449cc11, 32'hc2175ae0} /* (21, 21, 1) {real, imag} */,
  {32'hc4862669, 32'h00000000} /* (21, 21, 0) {real, imag} */,
  {32'h44a00c5f, 32'hc33a804c} /* (21, 20, 31) {real, imag} */,
  {32'hc4245fbb, 32'h42846104} /* (21, 20, 30) {real, imag} */,
  {32'hc2a03e4c, 32'h43276568} /* (21, 20, 29) {real, imag} */,
  {32'hc2ba0f3e, 32'hc2aabf02} /* (21, 20, 28) {real, imag} */,
  {32'hc2d8dcea, 32'h4284b96e} /* (21, 20, 27) {real, imag} */,
  {32'hc3020b5f, 32'hc3024399} /* (21, 20, 26) {real, imag} */,
  {32'h4233831a, 32'h420d953c} /* (21, 20, 25) {real, imag} */,
  {32'h42388039, 32'hc209b3cb} /* (21, 20, 24) {real, imag} */,
  {32'hc1c576ce, 32'h4282d49a} /* (21, 20, 23) {real, imag} */,
  {32'h4040ad78, 32'hc30e4bf0} /* (21, 20, 22) {real, imag} */,
  {32'h42291083, 32'h431cd1e4} /* (21, 20, 21) {real, imag} */,
  {32'h4197fcf8, 32'h41ce09ae} /* (21, 20, 20) {real, imag} */,
  {32'h41111380, 32'hc28abb72} /* (21, 20, 19) {real, imag} */,
  {32'h422b7d18, 32'hc27fbe00} /* (21, 20, 18) {real, imag} */,
  {32'hc2cace22, 32'hc21aa9f0} /* (21, 20, 17) {real, imag} */,
  {32'h428bdfdc, 32'h00000000} /* (21, 20, 16) {real, imag} */,
  {32'hc2cace22, 32'h421aa9f0} /* (21, 20, 15) {real, imag} */,
  {32'h422b7d18, 32'h427fbe00} /* (21, 20, 14) {real, imag} */,
  {32'h41111380, 32'h428abb72} /* (21, 20, 13) {real, imag} */,
  {32'h4197fcf8, 32'hc1ce09ae} /* (21, 20, 12) {real, imag} */,
  {32'h42291083, 32'hc31cd1e4} /* (21, 20, 11) {real, imag} */,
  {32'h4040ad78, 32'h430e4bf0} /* (21, 20, 10) {real, imag} */,
  {32'hc1c576ce, 32'hc282d49a} /* (21, 20, 9) {real, imag} */,
  {32'h42388039, 32'h4209b3cb} /* (21, 20, 8) {real, imag} */,
  {32'h4233831a, 32'hc20d953c} /* (21, 20, 7) {real, imag} */,
  {32'hc3020b5f, 32'h43024399} /* (21, 20, 6) {real, imag} */,
  {32'hc2d8dcea, 32'hc284b96e} /* (21, 20, 5) {real, imag} */,
  {32'hc2ba0f3e, 32'h42aabf02} /* (21, 20, 4) {real, imag} */,
  {32'hc2a03e4c, 32'hc3276568} /* (21, 20, 3) {real, imag} */,
  {32'hc4245fbb, 32'hc2846104} /* (21, 20, 2) {real, imag} */,
  {32'h44a00c5f, 32'h433a804c} /* (21, 20, 1) {real, imag} */,
  {32'h4392d1c4, 32'h00000000} /* (21, 20, 0) {real, imag} */,
  {32'h452a3934, 32'hc3f09bb4} /* (21, 19, 31) {real, imag} */,
  {32'hc488cf5e, 32'h43490f6c} /* (21, 19, 30) {real, imag} */,
  {32'h4062fbe0, 32'h425aa2b1} /* (21, 19, 29) {real, imag} */,
  {32'h427307fc, 32'hc21b379c} /* (21, 19, 28) {real, imag} */,
  {32'hc335bb87, 32'h42abece8} /* (21, 19, 27) {real, imag} */,
  {32'hc2bbcfca, 32'h41bc44fc} /* (21, 19, 26) {real, imag} */,
  {32'hc1c34476, 32'h42d38008} /* (21, 19, 25) {real, imag} */,
  {32'hc3184ac5, 32'h41a2238a} /* (21, 19, 24) {real, imag} */,
  {32'hc25dd2e1, 32'hc1c7035c} /* (21, 19, 23) {real, imag} */,
  {32'hc0d0709c, 32'hc2d79260} /* (21, 19, 22) {real, imag} */,
  {32'h41c63d5a, 32'hc1bdd0d6} /* (21, 19, 21) {real, imag} */,
  {32'h42b03115, 32'hc27397ac} /* (21, 19, 20) {real, imag} */,
  {32'hc28b42bf, 32'hc1dc2efc} /* (21, 19, 19) {real, imag} */,
  {32'hc0945098, 32'h41ccb82e} /* (21, 19, 18) {real, imag} */,
  {32'h41e11d90, 32'hc1ffc02d} /* (21, 19, 17) {real, imag} */,
  {32'h42223d52, 32'h00000000} /* (21, 19, 16) {real, imag} */,
  {32'h41e11d90, 32'h41ffc02d} /* (21, 19, 15) {real, imag} */,
  {32'hc0945098, 32'hc1ccb82e} /* (21, 19, 14) {real, imag} */,
  {32'hc28b42bf, 32'h41dc2efc} /* (21, 19, 13) {real, imag} */,
  {32'h42b03115, 32'h427397ac} /* (21, 19, 12) {real, imag} */,
  {32'h41c63d5a, 32'h41bdd0d6} /* (21, 19, 11) {real, imag} */,
  {32'hc0d0709c, 32'h42d79260} /* (21, 19, 10) {real, imag} */,
  {32'hc25dd2e1, 32'h41c7035c} /* (21, 19, 9) {real, imag} */,
  {32'hc3184ac5, 32'hc1a2238a} /* (21, 19, 8) {real, imag} */,
  {32'hc1c34476, 32'hc2d38008} /* (21, 19, 7) {real, imag} */,
  {32'hc2bbcfca, 32'hc1bc44fc} /* (21, 19, 6) {real, imag} */,
  {32'hc335bb87, 32'hc2abece8} /* (21, 19, 5) {real, imag} */,
  {32'h427307fc, 32'h421b379c} /* (21, 19, 4) {real, imag} */,
  {32'h4062fbe0, 32'hc25aa2b1} /* (21, 19, 3) {real, imag} */,
  {32'hc488cf5e, 32'hc3490f6c} /* (21, 19, 2) {real, imag} */,
  {32'h452a3934, 32'h43f09bb4} /* (21, 19, 1) {real, imag} */,
  {32'h449d0f4c, 32'h00000000} /* (21, 19, 0) {real, imag} */,
  {32'h45659d8b, 32'hc3f30184} /* (21, 18, 31) {real, imag} */,
  {32'hc4b13d7c, 32'h436ec7e5} /* (21, 18, 30) {real, imag} */,
  {32'h4086e3b0, 32'h42e82fc7} /* (21, 18, 29) {real, imag} */,
  {32'h42df42ca, 32'hc2ef717e} /* (21, 18, 28) {real, imag} */,
  {32'hc255de0a, 32'h42d01456} /* (21, 18, 27) {real, imag} */,
  {32'hc2c55101, 32'h42a0d55e} /* (21, 18, 26) {real, imag} */,
  {32'h42080322, 32'h42c8aaa5} /* (21, 18, 25) {real, imag} */,
  {32'hc1153340, 32'h42040dc4} /* (21, 18, 24) {real, imag} */,
  {32'hc263dc25, 32'hc070cee0} /* (21, 18, 23) {real, imag} */,
  {32'h417c3268, 32'h429911e9} /* (21, 18, 22) {real, imag} */,
  {32'hc21ee4ca, 32'hc34020f2} /* (21, 18, 21) {real, imag} */,
  {32'hc258eed0, 32'h428b51e6} /* (21, 18, 20) {real, imag} */,
  {32'h408b165a, 32'hc17fa339} /* (21, 18, 19) {real, imag} */,
  {32'hc1af1606, 32'hc2205bda} /* (21, 18, 18) {real, imag} */,
  {32'hc2618b59, 32'hc1ad794f} /* (21, 18, 17) {real, imag} */,
  {32'hc21a9c73, 32'h00000000} /* (21, 18, 16) {real, imag} */,
  {32'hc2618b59, 32'h41ad794f} /* (21, 18, 15) {real, imag} */,
  {32'hc1af1606, 32'h42205bda} /* (21, 18, 14) {real, imag} */,
  {32'h408b165a, 32'h417fa339} /* (21, 18, 13) {real, imag} */,
  {32'hc258eed0, 32'hc28b51e6} /* (21, 18, 12) {real, imag} */,
  {32'hc21ee4ca, 32'h434020f2} /* (21, 18, 11) {real, imag} */,
  {32'h417c3268, 32'hc29911e9} /* (21, 18, 10) {real, imag} */,
  {32'hc263dc25, 32'h4070cee0} /* (21, 18, 9) {real, imag} */,
  {32'hc1153340, 32'hc2040dc4} /* (21, 18, 8) {real, imag} */,
  {32'h42080322, 32'hc2c8aaa5} /* (21, 18, 7) {real, imag} */,
  {32'hc2c55101, 32'hc2a0d55e} /* (21, 18, 6) {real, imag} */,
  {32'hc255de0a, 32'hc2d01456} /* (21, 18, 5) {real, imag} */,
  {32'h42df42ca, 32'h42ef717e} /* (21, 18, 4) {real, imag} */,
  {32'h4086e3b0, 32'hc2e82fc7} /* (21, 18, 3) {real, imag} */,
  {32'hc4b13d7c, 32'hc36ec7e5} /* (21, 18, 2) {real, imag} */,
  {32'h45659d8b, 32'h43f30184} /* (21, 18, 1) {real, imag} */,
  {32'h450b3ad0, 32'h00000000} /* (21, 18, 0) {real, imag} */,
  {32'h458742d6, 32'hc4076aae} /* (21, 17, 31) {real, imag} */,
  {32'hc4c1a9f6, 32'h43a84092} /* (21, 17, 30) {real, imag} */,
  {32'hc1d96478, 32'h43913159} /* (21, 17, 29) {real, imag} */,
  {32'h4308d176, 32'hc30461aa} /* (21, 17, 28) {real, imag} */,
  {32'hc30f9474, 32'h436b872a} /* (21, 17, 27) {real, imag} */,
  {32'h41149c94, 32'h42264f72} /* (21, 17, 26) {real, imag} */,
  {32'h420d65ff, 32'h4326187f} /* (21, 17, 25) {real, imag} */,
  {32'h4231da78, 32'h42880235} /* (21, 17, 24) {real, imag} */,
  {32'hc2ab447f, 32'h42977de6} /* (21, 17, 23) {real, imag} */,
  {32'hc2905778, 32'h4214042c} /* (21, 17, 22) {real, imag} */,
  {32'hc22bd5a9, 32'h422f032a} /* (21, 17, 21) {real, imag} */,
  {32'hc16563ec, 32'hc266ac94} /* (21, 17, 20) {real, imag} */,
  {32'h4218538b, 32'h4182ecb8} /* (21, 17, 19) {real, imag} */,
  {32'h423ef4e1, 32'h42086004} /* (21, 17, 18) {real, imag} */,
  {32'hc293485e, 32'hc1cf0331} /* (21, 17, 17) {real, imag} */,
  {32'hc26b2c4e, 32'h00000000} /* (21, 17, 16) {real, imag} */,
  {32'hc293485e, 32'h41cf0331} /* (21, 17, 15) {real, imag} */,
  {32'h423ef4e1, 32'hc2086004} /* (21, 17, 14) {real, imag} */,
  {32'h4218538b, 32'hc182ecb8} /* (21, 17, 13) {real, imag} */,
  {32'hc16563ec, 32'h4266ac94} /* (21, 17, 12) {real, imag} */,
  {32'hc22bd5a9, 32'hc22f032a} /* (21, 17, 11) {real, imag} */,
  {32'hc2905778, 32'hc214042c} /* (21, 17, 10) {real, imag} */,
  {32'hc2ab447f, 32'hc2977de6} /* (21, 17, 9) {real, imag} */,
  {32'h4231da78, 32'hc2880235} /* (21, 17, 8) {real, imag} */,
  {32'h420d65ff, 32'hc326187f} /* (21, 17, 7) {real, imag} */,
  {32'h41149c94, 32'hc2264f72} /* (21, 17, 6) {real, imag} */,
  {32'hc30f9474, 32'hc36b872a} /* (21, 17, 5) {real, imag} */,
  {32'h4308d176, 32'h430461aa} /* (21, 17, 4) {real, imag} */,
  {32'hc1d96478, 32'hc3913159} /* (21, 17, 3) {real, imag} */,
  {32'hc4c1a9f6, 32'hc3a84092} /* (21, 17, 2) {real, imag} */,
  {32'h458742d6, 32'h44076aae} /* (21, 17, 1) {real, imag} */,
  {32'h452e1f78, 32'h00000000} /* (21, 17, 0) {real, imag} */,
  {32'h458df644, 32'hc3e09fb8} /* (21, 16, 31) {real, imag} */,
  {32'hc4bb78ba, 32'h43b74fe6} /* (21, 16, 30) {real, imag} */,
  {32'hc2d02b58, 32'h430561a4} /* (21, 16, 29) {real, imag} */,
  {32'h439ba107, 32'hc257bc85} /* (21, 16, 28) {real, imag} */,
  {32'hc3a2e972, 32'h423ca48e} /* (21, 16, 27) {real, imag} */,
  {32'h42e08d46, 32'h4252cb64} /* (21, 16, 26) {real, imag} */,
  {32'hc1f45928, 32'hc2226e04} /* (21, 16, 25) {real, imag} */,
  {32'hc1fec6bb, 32'h4306d587} /* (21, 16, 24) {real, imag} */,
  {32'hc29c2c15, 32'h424f4668} /* (21, 16, 23) {real, imag} */,
  {32'hc160a30d, 32'hc232c03a} /* (21, 16, 22) {real, imag} */,
  {32'h40491c70, 32'h428e7421} /* (21, 16, 21) {real, imag} */,
  {32'h42036c4b, 32'hc2649694} /* (21, 16, 20) {real, imag} */,
  {32'hc241ac1c, 32'h413cd702} /* (21, 16, 19) {real, imag} */,
  {32'h40d96b18, 32'h42d30eda} /* (21, 16, 18) {real, imag} */,
  {32'hc0e14900, 32'h42584c0a} /* (21, 16, 17) {real, imag} */,
  {32'h42421127, 32'h00000000} /* (21, 16, 16) {real, imag} */,
  {32'hc0e14900, 32'hc2584c0a} /* (21, 16, 15) {real, imag} */,
  {32'h40d96b18, 32'hc2d30eda} /* (21, 16, 14) {real, imag} */,
  {32'hc241ac1c, 32'hc13cd702} /* (21, 16, 13) {real, imag} */,
  {32'h42036c4b, 32'h42649694} /* (21, 16, 12) {real, imag} */,
  {32'h40491c70, 32'hc28e7421} /* (21, 16, 11) {real, imag} */,
  {32'hc160a30d, 32'h4232c03a} /* (21, 16, 10) {real, imag} */,
  {32'hc29c2c15, 32'hc24f4668} /* (21, 16, 9) {real, imag} */,
  {32'hc1fec6bb, 32'hc306d587} /* (21, 16, 8) {real, imag} */,
  {32'hc1f45928, 32'h42226e04} /* (21, 16, 7) {real, imag} */,
  {32'h42e08d46, 32'hc252cb64} /* (21, 16, 6) {real, imag} */,
  {32'hc3a2e972, 32'hc23ca48e} /* (21, 16, 5) {real, imag} */,
  {32'h439ba107, 32'h4257bc85} /* (21, 16, 4) {real, imag} */,
  {32'hc2d02b58, 32'hc30561a4} /* (21, 16, 3) {real, imag} */,
  {32'hc4bb78ba, 32'hc3b74fe6} /* (21, 16, 2) {real, imag} */,
  {32'h458df644, 32'h43e09fb8} /* (21, 16, 1) {real, imag} */,
  {32'h453dd41c, 32'h00000000} /* (21, 16, 0) {real, imag} */,
  {32'h458c83f8, 32'hc3def6a3} /* (21, 15, 31) {real, imag} */,
  {32'hc4b8fafa, 32'h43a2473a} /* (21, 15, 30) {real, imag} */,
  {32'hc31a74d4, 32'h42e3fb40} /* (21, 15, 29) {real, imag} */,
  {32'h43915360, 32'hc20051c8} /* (21, 15, 28) {real, imag} */,
  {32'hc38481ee, 32'h41eb8d30} /* (21, 15, 27) {real, imag} */,
  {32'hc22e7d67, 32'hc2e1879b} /* (21, 15, 26) {real, imag} */,
  {32'h41e3fcfb, 32'hc29b54b6} /* (21, 15, 25) {real, imag} */,
  {32'hc25628e0, 32'h42f842b7} /* (21, 15, 24) {real, imag} */,
  {32'h422dd25a, 32'h429bf45c} /* (21, 15, 23) {real, imag} */,
  {32'h42a2e3c8, 32'h41a13da9} /* (21, 15, 22) {real, imag} */,
  {32'hc2ec07c0, 32'h4254a8e6} /* (21, 15, 21) {real, imag} */,
  {32'hc2b5ca42, 32'h42aea814} /* (21, 15, 20) {real, imag} */,
  {32'hc2b35130, 32'h424fc49a} /* (21, 15, 19) {real, imag} */,
  {32'h420a7559, 32'h42cc45b6} /* (21, 15, 18) {real, imag} */,
  {32'h42000267, 32'hc295dcc8} /* (21, 15, 17) {real, imag} */,
  {32'hc2d04af9, 32'h00000000} /* (21, 15, 16) {real, imag} */,
  {32'h42000267, 32'h4295dcc8} /* (21, 15, 15) {real, imag} */,
  {32'h420a7559, 32'hc2cc45b6} /* (21, 15, 14) {real, imag} */,
  {32'hc2b35130, 32'hc24fc49a} /* (21, 15, 13) {real, imag} */,
  {32'hc2b5ca42, 32'hc2aea814} /* (21, 15, 12) {real, imag} */,
  {32'hc2ec07c0, 32'hc254a8e6} /* (21, 15, 11) {real, imag} */,
  {32'h42a2e3c8, 32'hc1a13da9} /* (21, 15, 10) {real, imag} */,
  {32'h422dd25a, 32'hc29bf45c} /* (21, 15, 9) {real, imag} */,
  {32'hc25628e0, 32'hc2f842b7} /* (21, 15, 8) {real, imag} */,
  {32'h41e3fcfb, 32'h429b54b6} /* (21, 15, 7) {real, imag} */,
  {32'hc22e7d67, 32'h42e1879b} /* (21, 15, 6) {real, imag} */,
  {32'hc38481ee, 32'hc1eb8d30} /* (21, 15, 5) {real, imag} */,
  {32'h43915360, 32'h420051c8} /* (21, 15, 4) {real, imag} */,
  {32'hc31a74d4, 32'hc2e3fb40} /* (21, 15, 3) {real, imag} */,
  {32'hc4b8fafa, 32'hc3a2473a} /* (21, 15, 2) {real, imag} */,
  {32'h458c83f8, 32'h43def6a3} /* (21, 15, 1) {real, imag} */,
  {32'h45443f04, 32'h00000000} /* (21, 15, 0) {real, imag} */,
  {32'h4583eb43, 32'hc3afa7cc} /* (21, 14, 31) {real, imag} */,
  {32'hc4b2f544, 32'h43adeee0} /* (21, 14, 30) {real, imag} */,
  {32'hc321ba46, 32'hc22a896a} /* (21, 14, 29) {real, imag} */,
  {32'h435f4beb, 32'hc2d06362} /* (21, 14, 28) {real, imag} */,
  {32'hc2e9a825, 32'h4343e649} /* (21, 14, 27) {real, imag} */,
  {32'hc2c3043b, 32'h405827c0} /* (21, 14, 26) {real, imag} */,
  {32'h419e2faf, 32'h40fa0c10} /* (21, 14, 25) {real, imag} */,
  {32'hc2965bc0, 32'h4341f98b} /* (21, 14, 24) {real, imag} */,
  {32'h416004fc, 32'h42f0d96b} /* (21, 14, 23) {real, imag} */,
  {32'hc221516c, 32'h424e16ae} /* (21, 14, 22) {real, imag} */,
  {32'hc2e57e93, 32'h42710196} /* (21, 14, 21) {real, imag} */,
  {32'hc06a7fa8, 32'hc20751e3} /* (21, 14, 20) {real, imag} */,
  {32'hc03f7e2c, 32'hc12f7d2d} /* (21, 14, 19) {real, imag} */,
  {32'h4234021d, 32'h410d37c6} /* (21, 14, 18) {real, imag} */,
  {32'hc27a5239, 32'hc233f338} /* (21, 14, 17) {real, imag} */,
  {32'hc16a0abb, 32'h00000000} /* (21, 14, 16) {real, imag} */,
  {32'hc27a5239, 32'h4233f338} /* (21, 14, 15) {real, imag} */,
  {32'h4234021d, 32'hc10d37c6} /* (21, 14, 14) {real, imag} */,
  {32'hc03f7e2c, 32'h412f7d2d} /* (21, 14, 13) {real, imag} */,
  {32'hc06a7fa8, 32'h420751e3} /* (21, 14, 12) {real, imag} */,
  {32'hc2e57e93, 32'hc2710196} /* (21, 14, 11) {real, imag} */,
  {32'hc221516c, 32'hc24e16ae} /* (21, 14, 10) {real, imag} */,
  {32'h416004fc, 32'hc2f0d96b} /* (21, 14, 9) {real, imag} */,
  {32'hc2965bc0, 32'hc341f98b} /* (21, 14, 8) {real, imag} */,
  {32'h419e2faf, 32'hc0fa0c10} /* (21, 14, 7) {real, imag} */,
  {32'hc2c3043b, 32'hc05827c0} /* (21, 14, 6) {real, imag} */,
  {32'hc2e9a825, 32'hc343e649} /* (21, 14, 5) {real, imag} */,
  {32'h435f4beb, 32'h42d06362} /* (21, 14, 4) {real, imag} */,
  {32'hc321ba46, 32'h422a896a} /* (21, 14, 3) {real, imag} */,
  {32'hc4b2f544, 32'hc3adeee0} /* (21, 14, 2) {real, imag} */,
  {32'h4583eb43, 32'h43afa7cc} /* (21, 14, 1) {real, imag} */,
  {32'h453e096c, 32'h00000000} /* (21, 14, 0) {real, imag} */,
  {32'h455c4a74, 32'hc32227f8} /* (21, 13, 31) {real, imag} */,
  {32'hc4acf42c, 32'h438c0d5c} /* (21, 13, 30) {real, imag} */,
  {32'hc2f49d88, 32'hc26a8d1b} /* (21, 13, 29) {real, imag} */,
  {32'h4393dace, 32'hc31c67c2} /* (21, 13, 28) {real, imag} */,
  {32'hc35b0e8d, 32'h438814bc} /* (21, 13, 27) {real, imag} */,
  {32'h429ceb22, 32'h42ce97e3} /* (21, 13, 26) {real, imag} */,
  {32'h42a80a24, 32'hc3101fde} /* (21, 13, 25) {real, imag} */,
  {32'hc1d4b408, 32'h42ed77d6} /* (21, 13, 24) {real, imag} */,
  {32'hc22633e1, 32'h430002e2} /* (21, 13, 23) {real, imag} */,
  {32'hc215d3d4, 32'h42c3139c} /* (21, 13, 22) {real, imag} */,
  {32'hc19a5efa, 32'h41a72ea2} /* (21, 13, 21) {real, imag} */,
  {32'hc18ad9d4, 32'h414bb518} /* (21, 13, 20) {real, imag} */,
  {32'h42fba83d, 32'hc247397a} /* (21, 13, 19) {real, imag} */,
  {32'hc2c88c52, 32'hc1b02a9e} /* (21, 13, 18) {real, imag} */,
  {32'hc283d1a5, 32'h422a59da} /* (21, 13, 17) {real, imag} */,
  {32'h42ae0cdb, 32'h00000000} /* (21, 13, 16) {real, imag} */,
  {32'hc283d1a5, 32'hc22a59da} /* (21, 13, 15) {real, imag} */,
  {32'hc2c88c52, 32'h41b02a9e} /* (21, 13, 14) {real, imag} */,
  {32'h42fba83d, 32'h4247397a} /* (21, 13, 13) {real, imag} */,
  {32'hc18ad9d4, 32'hc14bb518} /* (21, 13, 12) {real, imag} */,
  {32'hc19a5efa, 32'hc1a72ea2} /* (21, 13, 11) {real, imag} */,
  {32'hc215d3d4, 32'hc2c3139c} /* (21, 13, 10) {real, imag} */,
  {32'hc22633e1, 32'hc30002e2} /* (21, 13, 9) {real, imag} */,
  {32'hc1d4b408, 32'hc2ed77d6} /* (21, 13, 8) {real, imag} */,
  {32'h42a80a24, 32'h43101fde} /* (21, 13, 7) {real, imag} */,
  {32'h429ceb22, 32'hc2ce97e3} /* (21, 13, 6) {real, imag} */,
  {32'hc35b0e8d, 32'hc38814bc} /* (21, 13, 5) {real, imag} */,
  {32'h4393dace, 32'h431c67c2} /* (21, 13, 4) {real, imag} */,
  {32'hc2f49d88, 32'h426a8d1b} /* (21, 13, 3) {real, imag} */,
  {32'hc4acf42c, 32'hc38c0d5c} /* (21, 13, 2) {real, imag} */,
  {32'h455c4a74, 32'h432227f8} /* (21, 13, 1) {real, imag} */,
  {32'h45212bfe, 32'h00000000} /* (21, 13, 0) {real, imag} */,
  {32'h4516322a, 32'h42ddfdf8} /* (21, 12, 31) {real, imag} */,
  {32'hc4a02b56, 32'h431a2562} /* (21, 12, 30) {real, imag} */,
  {32'h42966f70, 32'hc1fd26f4} /* (21, 12, 29) {real, imag} */,
  {32'h437bee09, 32'hc2fd1eee} /* (21, 12, 28) {real, imag} */,
  {32'hc38e3018, 32'h42fcf446} /* (21, 12, 27) {real, imag} */,
  {32'h431ccc85, 32'h422329d4} /* (21, 12, 26) {real, imag} */,
  {32'h42e6fcb7, 32'hc2035440} /* (21, 12, 25) {real, imag} */,
  {32'h41fbac76, 32'hc1d9a826} /* (21, 12, 24) {real, imag} */,
  {32'hc2b102a4, 32'h429fa958} /* (21, 12, 23) {real, imag} */,
  {32'h4214dd68, 32'hc14f9358} /* (21, 12, 22) {real, imag} */,
  {32'hc2fa336a, 32'h43088000} /* (21, 12, 21) {real, imag} */,
  {32'hc25588ae, 32'h410e395c} /* (21, 12, 20) {real, imag} */,
  {32'h428d1ebd, 32'hc19b743a} /* (21, 12, 19) {real, imag} */,
  {32'hc27c1500, 32'h40d86350} /* (21, 12, 18) {real, imag} */,
  {32'h40afac10, 32'hc1ec5667} /* (21, 12, 17) {real, imag} */,
  {32'h3fdc6ea0, 32'h00000000} /* (21, 12, 16) {real, imag} */,
  {32'h40afac10, 32'h41ec5667} /* (21, 12, 15) {real, imag} */,
  {32'hc27c1500, 32'hc0d86350} /* (21, 12, 14) {real, imag} */,
  {32'h428d1ebd, 32'h419b743a} /* (21, 12, 13) {real, imag} */,
  {32'hc25588ae, 32'hc10e395c} /* (21, 12, 12) {real, imag} */,
  {32'hc2fa336a, 32'hc3088000} /* (21, 12, 11) {real, imag} */,
  {32'h4214dd68, 32'h414f9358} /* (21, 12, 10) {real, imag} */,
  {32'hc2b102a4, 32'hc29fa958} /* (21, 12, 9) {real, imag} */,
  {32'h41fbac76, 32'h41d9a826} /* (21, 12, 8) {real, imag} */,
  {32'h42e6fcb7, 32'h42035440} /* (21, 12, 7) {real, imag} */,
  {32'h431ccc85, 32'hc22329d4} /* (21, 12, 6) {real, imag} */,
  {32'hc38e3018, 32'hc2fcf446} /* (21, 12, 5) {real, imag} */,
  {32'h437bee09, 32'h42fd1eee} /* (21, 12, 4) {real, imag} */,
  {32'h42966f70, 32'h41fd26f4} /* (21, 12, 3) {real, imag} */,
  {32'hc4a02b56, 32'hc31a2562} /* (21, 12, 2) {real, imag} */,
  {32'h4516322a, 32'hc2ddfdf8} /* (21, 12, 1) {real, imag} */,
  {32'h44cfd0db, 32'h00000000} /* (21, 12, 0) {real, imag} */,
  {32'h448ba3c0, 32'h43f2d3e4} /* (21, 11, 31) {real, imag} */,
  {32'hc433bf26, 32'h4069b680} /* (21, 11, 30) {real, imag} */,
  {32'h425e8b76, 32'hc204a1ed} /* (21, 11, 29) {real, imag} */,
  {32'h4338ae39, 32'hc2e035a4} /* (21, 11, 28) {real, imag} */,
  {32'hc285fc80, 32'hc2223be3} /* (21, 11, 27) {real, imag} */,
  {32'h428119ef, 32'h4276e31a} /* (21, 11, 26) {real, imag} */,
  {32'h42461438, 32'h4229190a} /* (21, 11, 25) {real, imag} */,
  {32'hc303770d, 32'h42993211} /* (21, 11, 24) {real, imag} */,
  {32'h4025939c, 32'h41e7dcf8} /* (21, 11, 23) {real, imag} */,
  {32'h4285166a, 32'hc280bc29} /* (21, 11, 22) {real, imag} */,
  {32'hc30da14e, 32'h42a3a9db} /* (21, 11, 21) {real, imag} */,
  {32'hc28ebcff, 32'h421fed08} /* (21, 11, 20) {real, imag} */,
  {32'h42ba3854, 32'hc2457f95} /* (21, 11, 19) {real, imag} */,
  {32'hc2098e61, 32'hc1b9c84d} /* (21, 11, 18) {real, imag} */,
  {32'hc1b198b4, 32'h41c901ca} /* (21, 11, 17) {real, imag} */,
  {32'h428ead12, 32'h00000000} /* (21, 11, 16) {real, imag} */,
  {32'hc1b198b4, 32'hc1c901ca} /* (21, 11, 15) {real, imag} */,
  {32'hc2098e61, 32'h41b9c84d} /* (21, 11, 14) {real, imag} */,
  {32'h42ba3854, 32'h42457f95} /* (21, 11, 13) {real, imag} */,
  {32'hc28ebcff, 32'hc21fed08} /* (21, 11, 12) {real, imag} */,
  {32'hc30da14e, 32'hc2a3a9db} /* (21, 11, 11) {real, imag} */,
  {32'h4285166a, 32'h4280bc29} /* (21, 11, 10) {real, imag} */,
  {32'h4025939c, 32'hc1e7dcf8} /* (21, 11, 9) {real, imag} */,
  {32'hc303770d, 32'hc2993211} /* (21, 11, 8) {real, imag} */,
  {32'h42461438, 32'hc229190a} /* (21, 11, 7) {real, imag} */,
  {32'h428119ef, 32'hc276e31a} /* (21, 11, 6) {real, imag} */,
  {32'hc285fc80, 32'h42223be3} /* (21, 11, 5) {real, imag} */,
  {32'h4338ae39, 32'h42e035a4} /* (21, 11, 4) {real, imag} */,
  {32'h425e8b76, 32'h4204a1ed} /* (21, 11, 3) {real, imag} */,
  {32'hc433bf26, 32'hc069b680} /* (21, 11, 2) {real, imag} */,
  {32'h448ba3c0, 32'hc3f2d3e4} /* (21, 11, 1) {real, imag} */,
  {32'h44598ba2, 32'h00000000} /* (21, 11, 0) {real, imag} */,
  {32'hc42b7b08, 32'h444d888e} /* (21, 10, 31) {real, imag} */,
  {32'h431ac18c, 32'hc32c0cbc} /* (21, 10, 30) {real, imag} */,
  {32'h411bddf2, 32'hc195bea8} /* (21, 10, 29) {real, imag} */,
  {32'h4279bf3c, 32'hc27df095} /* (21, 10, 28) {real, imag} */,
  {32'h42fc9e82, 32'hc2819b9c} /* (21, 10, 27) {real, imag} */,
  {32'hc298eb1d, 32'h3fe612c0} /* (21, 10, 26) {real, imag} */,
  {32'hc31de222, 32'h42ac6f1c} /* (21, 10, 25) {real, imag} */,
  {32'h42368831, 32'hc28e2060} /* (21, 10, 24) {real, imag} */,
  {32'hc27f9a2e, 32'hc1c73b5f} /* (21, 10, 23) {real, imag} */,
  {32'hc10ecce6, 32'h41d0a34a} /* (21, 10, 22) {real, imag} */,
  {32'h417d7ad2, 32'hc2b93112} /* (21, 10, 21) {real, imag} */,
  {32'hc2b022cf, 32'hc25d82f4} /* (21, 10, 20) {real, imag} */,
  {32'hc217829e, 32'hc04facf2} /* (21, 10, 19) {real, imag} */,
  {32'h4214e448, 32'h41225e50} /* (21, 10, 18) {real, imag} */,
  {32'h41a74f9a, 32'hc1d7f507} /* (21, 10, 17) {real, imag} */,
  {32'h43019d02, 32'h00000000} /* (21, 10, 16) {real, imag} */,
  {32'h41a74f9a, 32'h41d7f507} /* (21, 10, 15) {real, imag} */,
  {32'h4214e448, 32'hc1225e50} /* (21, 10, 14) {real, imag} */,
  {32'hc217829e, 32'h404facf2} /* (21, 10, 13) {real, imag} */,
  {32'hc2b022cf, 32'h425d82f4} /* (21, 10, 12) {real, imag} */,
  {32'h417d7ad2, 32'h42b93112} /* (21, 10, 11) {real, imag} */,
  {32'hc10ecce6, 32'hc1d0a34a} /* (21, 10, 10) {real, imag} */,
  {32'hc27f9a2e, 32'h41c73b5f} /* (21, 10, 9) {real, imag} */,
  {32'h42368831, 32'h428e2060} /* (21, 10, 8) {real, imag} */,
  {32'hc31de222, 32'hc2ac6f1c} /* (21, 10, 7) {real, imag} */,
  {32'hc298eb1d, 32'hbfe612c0} /* (21, 10, 6) {real, imag} */,
  {32'h42fc9e82, 32'h42819b9c} /* (21, 10, 5) {real, imag} */,
  {32'h4279bf3c, 32'h427df095} /* (21, 10, 4) {real, imag} */,
  {32'h411bddf2, 32'h4195bea8} /* (21, 10, 3) {real, imag} */,
  {32'h431ac18c, 32'h432c0cbc} /* (21, 10, 2) {real, imag} */,
  {32'hc42b7b08, 32'hc44d888e} /* (21, 10, 1) {real, imag} */,
  {32'hc453598d, 32'h00000000} /* (21, 10, 0) {real, imag} */,
  {32'hc508dd34, 32'h44829d78} /* (21, 9, 31) {real, imag} */,
  {32'h444794c2, 32'hc3be49e0} /* (21, 9, 30) {real, imag} */,
  {32'h42d4b6a6, 32'hbe384740} /* (21, 9, 29) {real, imag} */,
  {32'h3f673000, 32'h42e0e58a} /* (21, 9, 28) {real, imag} */,
  {32'h431ad770, 32'hc2247cf3} /* (21, 9, 27) {real, imag} */,
  {32'h4274c9d0, 32'hc29a57e2} /* (21, 9, 26) {real, imag} */,
  {32'hc2aaf224, 32'h42eae69c} /* (21, 9, 25) {real, imag} */,
  {32'h429dd0a6, 32'hc2ef4344} /* (21, 9, 24) {real, imag} */,
  {32'hc28b1c76, 32'hc25937cc} /* (21, 9, 23) {real, imag} */,
  {32'hc1a02f1e, 32'h4223d408} /* (21, 9, 22) {real, imag} */,
  {32'hc2e1c88f, 32'hc29bf294} /* (21, 9, 21) {real, imag} */,
  {32'h4095a7ca, 32'h423926e4} /* (21, 9, 20) {real, imag} */,
  {32'h426bd6f8, 32'h42ad1369} /* (21, 9, 19) {real, imag} */,
  {32'h3e8284a0, 32'h420e2e12} /* (21, 9, 18) {real, imag} */,
  {32'hc26161ca, 32'h42e6de0b} /* (21, 9, 17) {real, imag} */,
  {32'h421dc04a, 32'h00000000} /* (21, 9, 16) {real, imag} */,
  {32'hc26161ca, 32'hc2e6de0b} /* (21, 9, 15) {real, imag} */,
  {32'h3e8284a0, 32'hc20e2e12} /* (21, 9, 14) {real, imag} */,
  {32'h426bd6f8, 32'hc2ad1369} /* (21, 9, 13) {real, imag} */,
  {32'h4095a7ca, 32'hc23926e4} /* (21, 9, 12) {real, imag} */,
  {32'hc2e1c88f, 32'h429bf294} /* (21, 9, 11) {real, imag} */,
  {32'hc1a02f1e, 32'hc223d408} /* (21, 9, 10) {real, imag} */,
  {32'hc28b1c76, 32'h425937cc} /* (21, 9, 9) {real, imag} */,
  {32'h429dd0a6, 32'h42ef4344} /* (21, 9, 8) {real, imag} */,
  {32'hc2aaf224, 32'hc2eae69c} /* (21, 9, 7) {real, imag} */,
  {32'h4274c9d0, 32'h429a57e2} /* (21, 9, 6) {real, imag} */,
  {32'h431ad770, 32'h42247cf3} /* (21, 9, 5) {real, imag} */,
  {32'h3f673000, 32'hc2e0e58a} /* (21, 9, 4) {real, imag} */,
  {32'h42d4b6a6, 32'h3e384740} /* (21, 9, 3) {real, imag} */,
  {32'h444794c2, 32'h43be49e0} /* (21, 9, 2) {real, imag} */,
  {32'hc508dd34, 32'hc4829d78} /* (21, 9, 1) {real, imag} */,
  {32'hc5120600, 32'h00000000} /* (21, 9, 0) {real, imag} */,
  {32'hc543a334, 32'h44c99c3f} /* (21, 8, 31) {real, imag} */,
  {32'h44763c20, 32'hc3dc0184} /* (21, 8, 30) {real, imag} */,
  {32'h3efc6f00, 32'hc10ee248} /* (21, 8, 29) {real, imag} */,
  {32'h40f9e030, 32'h430daf44} /* (21, 8, 28) {real, imag} */,
  {32'h4353707c, 32'hc2e0095a} /* (21, 8, 27) {real, imag} */,
  {32'h4254343b, 32'hc2949cea} /* (21, 8, 26) {real, imag} */,
  {32'h425fd8a0, 32'h4282cf5a} /* (21, 8, 25) {real, imag} */,
  {32'h42785540, 32'hc34315d6} /* (21, 8, 24) {real, imag} */,
  {32'h42801cb0, 32'hc031a840} /* (21, 8, 23) {real, imag} */,
  {32'hc1b7947c, 32'h42df2ecf} /* (21, 8, 22) {real, imag} */,
  {32'h42530d72, 32'hc08ab524} /* (21, 8, 21) {real, imag} */,
  {32'h419acc70, 32'h421ebf94} /* (21, 8, 20) {real, imag} */,
  {32'h423aa243, 32'hc1dfba44} /* (21, 8, 19) {real, imag} */,
  {32'hc1df15ac, 32'hc25c0b15} /* (21, 8, 18) {real, imag} */,
  {32'h42a1dc0c, 32'h4236f1b5} /* (21, 8, 17) {real, imag} */,
  {32'hc204586f, 32'h00000000} /* (21, 8, 16) {real, imag} */,
  {32'h42a1dc0c, 32'hc236f1b5} /* (21, 8, 15) {real, imag} */,
  {32'hc1df15ac, 32'h425c0b15} /* (21, 8, 14) {real, imag} */,
  {32'h423aa243, 32'h41dfba44} /* (21, 8, 13) {real, imag} */,
  {32'h419acc70, 32'hc21ebf94} /* (21, 8, 12) {real, imag} */,
  {32'h42530d72, 32'h408ab524} /* (21, 8, 11) {real, imag} */,
  {32'hc1b7947c, 32'hc2df2ecf} /* (21, 8, 10) {real, imag} */,
  {32'h42801cb0, 32'h4031a840} /* (21, 8, 9) {real, imag} */,
  {32'h42785540, 32'h434315d6} /* (21, 8, 8) {real, imag} */,
  {32'h425fd8a0, 32'hc282cf5a} /* (21, 8, 7) {real, imag} */,
  {32'h4254343b, 32'h42949cea} /* (21, 8, 6) {real, imag} */,
  {32'h4353707c, 32'h42e0095a} /* (21, 8, 5) {real, imag} */,
  {32'h40f9e030, 32'hc30daf44} /* (21, 8, 4) {real, imag} */,
  {32'h3efc6f00, 32'h410ee248} /* (21, 8, 3) {real, imag} */,
  {32'h44763c20, 32'h43dc0184} /* (21, 8, 2) {real, imag} */,
  {32'hc543a334, 32'hc4c99c3f} /* (21, 8, 1) {real, imag} */,
  {32'hc54622dc, 32'h00000000} /* (21, 8, 0) {real, imag} */,
  {32'hc56d0d36, 32'h4501c2b2} /* (21, 7, 31) {real, imag} */,
  {32'h44745fb4, 32'hc40b5481} /* (21, 7, 30) {real, imag} */,
  {32'h409a4008, 32'hc20d6621} /* (21, 7, 29) {real, imag} */,
  {32'hc1678d80, 32'h4248b68a} /* (21, 7, 28) {real, imag} */,
  {32'h431adf34, 32'h41e48fa4} /* (21, 7, 27) {real, imag} */,
  {32'h41a429d7, 32'h417efe24} /* (21, 7, 26) {real, imag} */,
  {32'h42d14ab7, 32'h4235c01e} /* (21, 7, 25) {real, imag} */,
  {32'h42b60a26, 32'hc3238f41} /* (21, 7, 24) {real, imag} */,
  {32'hc0ffc658, 32'hc26d988c} /* (21, 7, 23) {real, imag} */,
  {32'h420ccb1f, 32'hc22c27c0} /* (21, 7, 22) {real, imag} */,
  {32'h41514f90, 32'h414425d4} /* (21, 7, 21) {real, imag} */,
  {32'hc1233b08, 32'h40a3aa40} /* (21, 7, 20) {real, imag} */,
  {32'h40d29acc, 32'h424b00a5} /* (21, 7, 19) {real, imag} */,
  {32'h4278d97f, 32'h423958ce} /* (21, 7, 18) {real, imag} */,
  {32'hc26e8f09, 32'h4195a63c} /* (21, 7, 17) {real, imag} */,
  {32'h42ad2248, 32'h00000000} /* (21, 7, 16) {real, imag} */,
  {32'hc26e8f09, 32'hc195a63c} /* (21, 7, 15) {real, imag} */,
  {32'h4278d97f, 32'hc23958ce} /* (21, 7, 14) {real, imag} */,
  {32'h40d29acc, 32'hc24b00a5} /* (21, 7, 13) {real, imag} */,
  {32'hc1233b08, 32'hc0a3aa40} /* (21, 7, 12) {real, imag} */,
  {32'h41514f90, 32'hc14425d4} /* (21, 7, 11) {real, imag} */,
  {32'h420ccb1f, 32'h422c27c0} /* (21, 7, 10) {real, imag} */,
  {32'hc0ffc658, 32'h426d988c} /* (21, 7, 9) {real, imag} */,
  {32'h42b60a26, 32'h43238f41} /* (21, 7, 8) {real, imag} */,
  {32'h42d14ab7, 32'hc235c01e} /* (21, 7, 7) {real, imag} */,
  {32'h41a429d7, 32'hc17efe24} /* (21, 7, 6) {real, imag} */,
  {32'h431adf34, 32'hc1e48fa4} /* (21, 7, 5) {real, imag} */,
  {32'hc1678d80, 32'hc248b68a} /* (21, 7, 4) {real, imag} */,
  {32'h409a4008, 32'h420d6621} /* (21, 7, 3) {real, imag} */,
  {32'h44745fb4, 32'h440b5481} /* (21, 7, 2) {real, imag} */,
  {32'hc56d0d36, 32'hc501c2b2} /* (21, 7, 1) {real, imag} */,
  {32'hc57ca1ee, 32'h00000000} /* (21, 7, 0) {real, imag} */,
  {32'hc578d328, 32'h451b5521} /* (21, 6, 31) {real, imag} */,
  {32'h445fa9e1, 32'hc43594bc} /* (21, 6, 30) {real, imag} */,
  {32'hc1b52e29, 32'hc28b837f} /* (21, 6, 29) {real, imag} */,
  {32'hc1a520f0, 32'hc32fc0f2} /* (21, 6, 28) {real, imag} */,
  {32'h4330a375, 32'hc2031fdc} /* (21, 6, 27) {real, imag} */,
  {32'hc2a8de43, 32'h3fdc24f0} /* (21, 6, 26) {real, imag} */,
  {32'h42df826b, 32'h41cda744} /* (21, 6, 25) {real, imag} */,
  {32'h4102546c, 32'hc20e3cb0} /* (21, 6, 24) {real, imag} */,
  {32'h424159f2, 32'h424d5fca} /* (21, 6, 23) {real, imag} */,
  {32'h42918206, 32'h430311e2} /* (21, 6, 22) {real, imag} */,
  {32'hc16dc84c, 32'h4294edf3} /* (21, 6, 21) {real, imag} */,
  {32'hc23fc808, 32'hc2af3426} /* (21, 6, 20) {real, imag} */,
  {32'hc125c5f7, 32'h40e49cc4} /* (21, 6, 19) {real, imag} */,
  {32'h41482ed0, 32'hc27730a0} /* (21, 6, 18) {real, imag} */,
  {32'h41cfc683, 32'h42ab5562} /* (21, 6, 17) {real, imag} */,
  {32'hc07df608, 32'h00000000} /* (21, 6, 16) {real, imag} */,
  {32'h41cfc683, 32'hc2ab5562} /* (21, 6, 15) {real, imag} */,
  {32'h41482ed0, 32'h427730a0} /* (21, 6, 14) {real, imag} */,
  {32'hc125c5f7, 32'hc0e49cc4} /* (21, 6, 13) {real, imag} */,
  {32'hc23fc808, 32'h42af3426} /* (21, 6, 12) {real, imag} */,
  {32'hc16dc84c, 32'hc294edf3} /* (21, 6, 11) {real, imag} */,
  {32'h42918206, 32'hc30311e2} /* (21, 6, 10) {real, imag} */,
  {32'h424159f2, 32'hc24d5fca} /* (21, 6, 9) {real, imag} */,
  {32'h4102546c, 32'h420e3cb0} /* (21, 6, 8) {real, imag} */,
  {32'h42df826b, 32'hc1cda744} /* (21, 6, 7) {real, imag} */,
  {32'hc2a8de43, 32'hbfdc24f0} /* (21, 6, 6) {real, imag} */,
  {32'h4330a375, 32'h42031fdc} /* (21, 6, 5) {real, imag} */,
  {32'hc1a520f0, 32'h432fc0f2} /* (21, 6, 4) {real, imag} */,
  {32'hc1b52e29, 32'h428b837f} /* (21, 6, 3) {real, imag} */,
  {32'h445fa9e1, 32'h443594bc} /* (21, 6, 2) {real, imag} */,
  {32'hc578d328, 32'hc51b5521} /* (21, 6, 1) {real, imag} */,
  {32'hc589d7f9, 32'h00000000} /* (21, 6, 0) {real, imag} */,
  {32'hc573ca9b, 32'h45525d84} /* (21, 5, 31) {real, imag} */,
  {32'h438b6638, 32'hc467149b} /* (21, 5, 30) {real, imag} */,
  {32'h42824b19, 32'hc30b0598} /* (21, 5, 29) {real, imag} */,
  {32'h434566fe, 32'hc349954d} /* (21, 5, 28) {real, imag} */,
  {32'h43364c48, 32'h425f2c92} /* (21, 5, 27) {real, imag} */,
  {32'hc303d81d, 32'h4283fd22} /* (21, 5, 26) {real, imag} */,
  {32'h42bb7793, 32'h4296d138} /* (21, 5, 25) {real, imag} */,
  {32'hc0caf9f4, 32'hc2fa352e} /* (21, 5, 24) {real, imag} */,
  {32'h421dedf3, 32'h41f64eb4} /* (21, 5, 23) {real, imag} */,
  {32'hc1ad34d2, 32'h413f0654} /* (21, 5, 22) {real, imag} */,
  {32'hc2cc5b91, 32'hc21d90f4} /* (21, 5, 21) {real, imag} */,
  {32'hc067f3c0, 32'hc29f186a} /* (21, 5, 20) {real, imag} */,
  {32'h4213ef41, 32'h41d04104} /* (21, 5, 19) {real, imag} */,
  {32'hc0de88b0, 32'hc1895cbc} /* (21, 5, 18) {real, imag} */,
  {32'hc15bd6c5, 32'h41d0599f} /* (21, 5, 17) {real, imag} */,
  {32'h4119ec80, 32'h00000000} /* (21, 5, 16) {real, imag} */,
  {32'hc15bd6c5, 32'hc1d0599f} /* (21, 5, 15) {real, imag} */,
  {32'hc0de88b0, 32'h41895cbc} /* (21, 5, 14) {real, imag} */,
  {32'h4213ef41, 32'hc1d04104} /* (21, 5, 13) {real, imag} */,
  {32'hc067f3c0, 32'h429f186a} /* (21, 5, 12) {real, imag} */,
  {32'hc2cc5b91, 32'h421d90f4} /* (21, 5, 11) {real, imag} */,
  {32'hc1ad34d2, 32'hc13f0654} /* (21, 5, 10) {real, imag} */,
  {32'h421dedf3, 32'hc1f64eb4} /* (21, 5, 9) {real, imag} */,
  {32'hc0caf9f4, 32'h42fa352e} /* (21, 5, 8) {real, imag} */,
  {32'h42bb7793, 32'hc296d138} /* (21, 5, 7) {real, imag} */,
  {32'hc303d81d, 32'hc283fd22} /* (21, 5, 6) {real, imag} */,
  {32'h43364c48, 32'hc25f2c92} /* (21, 5, 5) {real, imag} */,
  {32'h434566fe, 32'h4349954d} /* (21, 5, 4) {real, imag} */,
  {32'h42824b19, 32'h430b0598} /* (21, 5, 3) {real, imag} */,
  {32'h438b6638, 32'h4467149b} /* (21, 5, 2) {real, imag} */,
  {32'hc573ca9b, 32'hc5525d84} /* (21, 5, 1) {real, imag} */,
  {32'hc5955c8b, 32'h00000000} /* (21, 5, 0) {real, imag} */,
  {32'hc55f0c5c, 32'h45749b6d} /* (21, 4, 31) {real, imag} */,
  {32'hc2bec1c8, 32'hc4886e2d} /* (21, 4, 30) {real, imag} */,
  {32'h42ecd48c, 32'hc3531bc0} /* (21, 4, 29) {real, imag} */,
  {32'h42d633fa, 32'hc3dddd09} /* (21, 4, 28) {real, imag} */,
  {32'h42c1b2ac, 32'h4276aac8} /* (21, 4, 27) {real, imag} */,
  {32'h42a65b7a, 32'h4259af8d} /* (21, 4, 26) {real, imag} */,
  {32'h42dbd7c6, 32'hc1597644} /* (21, 4, 25) {real, imag} */,
  {32'hc3214392, 32'h41e45396} /* (21, 4, 24) {real, imag} */,
  {32'h42f71414, 32'hc247701c} /* (21, 4, 23) {real, imag} */,
  {32'h42503f89, 32'h41985670} /* (21, 4, 22) {real, imag} */,
  {32'hc2b17c22, 32'h41d954ba} /* (21, 4, 21) {real, imag} */,
  {32'hc2bfea43, 32'h429364b5} /* (21, 4, 20) {real, imag} */,
  {32'hc099ccf8, 32'hc0443030} /* (21, 4, 19) {real, imag} */,
  {32'hc14ce940, 32'hc069a564} /* (21, 4, 18) {real, imag} */,
  {32'hc0ccd8a0, 32'hc20b26ba} /* (21, 4, 17) {real, imag} */,
  {32'hc1a45942, 32'h00000000} /* (21, 4, 16) {real, imag} */,
  {32'hc0ccd8a0, 32'h420b26ba} /* (21, 4, 15) {real, imag} */,
  {32'hc14ce940, 32'h4069a564} /* (21, 4, 14) {real, imag} */,
  {32'hc099ccf8, 32'h40443030} /* (21, 4, 13) {real, imag} */,
  {32'hc2bfea43, 32'hc29364b5} /* (21, 4, 12) {real, imag} */,
  {32'hc2b17c22, 32'hc1d954ba} /* (21, 4, 11) {real, imag} */,
  {32'h42503f89, 32'hc1985670} /* (21, 4, 10) {real, imag} */,
  {32'h42f71414, 32'h4247701c} /* (21, 4, 9) {real, imag} */,
  {32'hc3214392, 32'hc1e45396} /* (21, 4, 8) {real, imag} */,
  {32'h42dbd7c6, 32'h41597644} /* (21, 4, 7) {real, imag} */,
  {32'h42a65b7a, 32'hc259af8d} /* (21, 4, 6) {real, imag} */,
  {32'h42c1b2ac, 32'hc276aac8} /* (21, 4, 5) {real, imag} */,
  {32'h42d633fa, 32'h43dddd09} /* (21, 4, 4) {real, imag} */,
  {32'h42ecd48c, 32'h43531bc0} /* (21, 4, 3) {real, imag} */,
  {32'hc2bec1c8, 32'h44886e2d} /* (21, 4, 2) {real, imag} */,
  {32'hc55f0c5c, 32'hc5749b6d} /* (21, 4, 1) {real, imag} */,
  {32'hc5a4c735, 32'h00000000} /* (21, 4, 0) {real, imag} */,
  {32'hc55f470e, 32'h4580f8e8} /* (21, 3, 31) {real, imag} */,
  {32'hc3a63174, 32'hc481e7fa} /* (21, 3, 30) {real, imag} */,
  {32'h41111498, 32'hc2c12c13} /* (21, 3, 29) {real, imag} */,
  {32'h4298c176, 32'hc3cba501} /* (21, 3, 28) {real, imag} */,
  {32'h43a12b3e, 32'h42f8958c} /* (21, 3, 27) {real, imag} */,
  {32'h419e9359, 32'hc28368e8} /* (21, 3, 26) {real, imag} */,
  {32'h4129f10b, 32'h426e7201} /* (21, 3, 25) {real, imag} */,
  {32'hc1bc0ecb, 32'hc2bc427e} /* (21, 3, 24) {real, imag} */,
  {32'h430c2208, 32'h421a998d} /* (21, 3, 23) {real, imag} */,
  {32'h4292ddd3, 32'hc1e18a78} /* (21, 3, 22) {real, imag} */,
  {32'h41f4ee34, 32'hc1daf740} /* (21, 3, 21) {real, imag} */,
  {32'hc2552e86, 32'hc2e865fd} /* (21, 3, 20) {real, imag} */,
  {32'h41465026, 32'hc25b95e3} /* (21, 3, 19) {real, imag} */,
  {32'h4283e030, 32'hc2bdf4e4} /* (21, 3, 18) {real, imag} */,
  {32'h410bf682, 32'h41704dcc} /* (21, 3, 17) {real, imag} */,
  {32'h41982cbb, 32'h00000000} /* (21, 3, 16) {real, imag} */,
  {32'h410bf682, 32'hc1704dcc} /* (21, 3, 15) {real, imag} */,
  {32'h4283e030, 32'h42bdf4e4} /* (21, 3, 14) {real, imag} */,
  {32'h41465026, 32'h425b95e3} /* (21, 3, 13) {real, imag} */,
  {32'hc2552e86, 32'h42e865fd} /* (21, 3, 12) {real, imag} */,
  {32'h41f4ee34, 32'h41daf740} /* (21, 3, 11) {real, imag} */,
  {32'h4292ddd3, 32'h41e18a78} /* (21, 3, 10) {real, imag} */,
  {32'h430c2208, 32'hc21a998d} /* (21, 3, 9) {real, imag} */,
  {32'hc1bc0ecb, 32'h42bc427e} /* (21, 3, 8) {real, imag} */,
  {32'h4129f10b, 32'hc26e7201} /* (21, 3, 7) {real, imag} */,
  {32'h419e9359, 32'h428368e8} /* (21, 3, 6) {real, imag} */,
  {32'h43a12b3e, 32'hc2f8958c} /* (21, 3, 5) {real, imag} */,
  {32'h4298c176, 32'h43cba501} /* (21, 3, 4) {real, imag} */,
  {32'h41111498, 32'h42c12c13} /* (21, 3, 3) {real, imag} */,
  {32'hc3a63174, 32'h4481e7fa} /* (21, 3, 2) {real, imag} */,
  {32'hc55f470e, 32'hc580f8e8} /* (21, 3, 1) {real, imag} */,
  {32'hc5ae27c6, 32'h00000000} /* (21, 3, 0) {real, imag} */,
  {32'hc55ea37c, 32'h457a541a} /* (21, 2, 31) {real, imag} */,
  {32'hc38a4e0a, 32'hc475b01e} /* (21, 2, 30) {real, imag} */,
  {32'h41816884, 32'hc3293158} /* (21, 2, 29) {real, imag} */,
  {32'h42dc4a03, 32'hc38a40c2} /* (21, 2, 28) {real, imag} */,
  {32'h4367f41b, 32'h4267951a} /* (21, 2, 27) {real, imag} */,
  {32'h42029a62, 32'hc17b0748} /* (21, 2, 26) {real, imag} */,
  {32'h42c854f8, 32'hc13c4cfe} /* (21, 2, 25) {real, imag} */,
  {32'hc1e923cb, 32'hc283b4fa} /* (21, 2, 24) {real, imag} */,
  {32'h41a0c256, 32'hc27d0c4e} /* (21, 2, 23) {real, imag} */,
  {32'h427d5037, 32'hc113b800} /* (21, 2, 22) {real, imag} */,
  {32'h42c3083e, 32'hc21d0d67} /* (21, 2, 21) {real, imag} */,
  {32'h4210c77c, 32'h41ac7390} /* (21, 2, 20) {real, imag} */,
  {32'h42706eba, 32'h41a63322} /* (21, 2, 19) {real, imag} */,
  {32'hc184f474, 32'h40e22bbc} /* (21, 2, 18) {real, imag} */,
  {32'hc15ed70c, 32'h42828ea9} /* (21, 2, 17) {real, imag} */,
  {32'h3e88f600, 32'h00000000} /* (21, 2, 16) {real, imag} */,
  {32'hc15ed70c, 32'hc2828ea9} /* (21, 2, 15) {real, imag} */,
  {32'hc184f474, 32'hc0e22bbc} /* (21, 2, 14) {real, imag} */,
  {32'h42706eba, 32'hc1a63322} /* (21, 2, 13) {real, imag} */,
  {32'h4210c77c, 32'hc1ac7390} /* (21, 2, 12) {real, imag} */,
  {32'h42c3083e, 32'h421d0d67} /* (21, 2, 11) {real, imag} */,
  {32'h427d5037, 32'h4113b800} /* (21, 2, 10) {real, imag} */,
  {32'h41a0c256, 32'h427d0c4e} /* (21, 2, 9) {real, imag} */,
  {32'hc1e923cb, 32'h4283b4fa} /* (21, 2, 8) {real, imag} */,
  {32'h42c854f8, 32'h413c4cfe} /* (21, 2, 7) {real, imag} */,
  {32'h42029a62, 32'h417b0748} /* (21, 2, 6) {real, imag} */,
  {32'h4367f41b, 32'hc267951a} /* (21, 2, 5) {real, imag} */,
  {32'h42dc4a03, 32'h438a40c2} /* (21, 2, 4) {real, imag} */,
  {32'h41816884, 32'h43293158} /* (21, 2, 3) {real, imag} */,
  {32'hc38a4e0a, 32'h4475b01e} /* (21, 2, 2) {real, imag} */,
  {32'hc55ea37c, 32'hc57a541a} /* (21, 2, 1) {real, imag} */,
  {32'hc5ae2d8e, 32'h00000000} /* (21, 2, 0) {real, imag} */,
  {32'hc5631050, 32'h456ec5da} /* (21, 1, 31) {real, imag} */,
  {32'h40c79180, 32'hc470b41f} /* (21, 1, 30) {real, imag} */,
  {32'h431a3542, 32'hc30163f5} /* (21, 1, 29) {real, imag} */,
  {32'h42de13e9, 32'hc3693a30} /* (21, 1, 28) {real, imag} */,
  {32'h4380d744, 32'hc251db61} /* (21, 1, 27) {real, imag} */,
  {32'h4291a8c3, 32'hc28aa9d3} /* (21, 1, 26) {real, imag} */,
  {32'h42bca11f, 32'h41686b7c} /* (21, 1, 25) {real, imag} */,
  {32'hc28d2ba7, 32'h4242a8fe} /* (21, 1, 24) {real, imag} */,
  {32'h421d879a, 32'hc1d209b6} /* (21, 1, 23) {real, imag} */,
  {32'hc0368e0e, 32'hc23db598} /* (21, 1, 22) {real, imag} */,
  {32'h41b2f558, 32'h424228da} /* (21, 1, 21) {real, imag} */,
  {32'hc1f7480f, 32'h42ca7983} /* (21, 1, 20) {real, imag} */,
  {32'h41bdfc3b, 32'h418b346e} /* (21, 1, 19) {real, imag} */,
  {32'hc29d6379, 32'h4286f9a4} /* (21, 1, 18) {real, imag} */,
  {32'h41aa645e, 32'hc22c72fa} /* (21, 1, 17) {real, imag} */,
  {32'h42a78712, 32'h00000000} /* (21, 1, 16) {real, imag} */,
  {32'h41aa645e, 32'h422c72fa} /* (21, 1, 15) {real, imag} */,
  {32'hc29d6379, 32'hc286f9a4} /* (21, 1, 14) {real, imag} */,
  {32'h41bdfc3b, 32'hc18b346e} /* (21, 1, 13) {real, imag} */,
  {32'hc1f7480f, 32'hc2ca7983} /* (21, 1, 12) {real, imag} */,
  {32'h41b2f558, 32'hc24228da} /* (21, 1, 11) {real, imag} */,
  {32'hc0368e0e, 32'h423db598} /* (21, 1, 10) {real, imag} */,
  {32'h421d879a, 32'h41d209b6} /* (21, 1, 9) {real, imag} */,
  {32'hc28d2ba7, 32'hc242a8fe} /* (21, 1, 8) {real, imag} */,
  {32'h42bca11f, 32'hc1686b7c} /* (21, 1, 7) {real, imag} */,
  {32'h4291a8c3, 32'h428aa9d3} /* (21, 1, 6) {real, imag} */,
  {32'h4380d744, 32'h4251db61} /* (21, 1, 5) {real, imag} */,
  {32'h42de13e9, 32'h43693a30} /* (21, 1, 4) {real, imag} */,
  {32'h431a3542, 32'h430163f5} /* (21, 1, 3) {real, imag} */,
  {32'h40c79180, 32'h4470b41f} /* (21, 1, 2) {real, imag} */,
  {32'hc5631050, 32'hc56ec5da} /* (21, 1, 1) {real, imag} */,
  {32'hc5b1b29b, 32'h00000000} /* (21, 1, 0) {real, imag} */,
  {32'hc56c4589, 32'h4545a4e8} /* (21, 0, 31) {real, imag} */,
  {32'h4380d046, 32'hc4430249} /* (21, 0, 30) {real, imag} */,
  {32'h43619e64, 32'h419b2a64} /* (21, 0, 29) {real, imag} */,
  {32'hc18babf0, 32'hc32716b9} /* (21, 0, 28) {real, imag} */,
  {32'h42a63412, 32'hc1e3c34c} /* (21, 0, 27) {real, imag} */,
  {32'hc2745329, 32'hc1dc03bc} /* (21, 0, 26) {real, imag} */,
  {32'hc1aa5fd4, 32'h42af723a} /* (21, 0, 25) {real, imag} */,
  {32'hc1c182df, 32'h3fee5680} /* (21, 0, 24) {real, imag} */,
  {32'h4289386d, 32'hc0a366ac} /* (21, 0, 23) {real, imag} */,
  {32'h417a010b, 32'hc31d13b6} /* (21, 0, 22) {real, imag} */,
  {32'hc2144a57, 32'h42722322} /* (21, 0, 21) {real, imag} */,
  {32'h423f9fc9, 32'hc27f0f22} /* (21, 0, 20) {real, imag} */,
  {32'hc13b46ba, 32'h41d0075f} /* (21, 0, 19) {real, imag} */,
  {32'h4216714d, 32'h40fb7bd0} /* (21, 0, 18) {real, imag} */,
  {32'h41cc1b98, 32'h41af4617} /* (21, 0, 17) {real, imag} */,
  {32'hc280305f, 32'h00000000} /* (21, 0, 16) {real, imag} */,
  {32'h41cc1b98, 32'hc1af4617} /* (21, 0, 15) {real, imag} */,
  {32'h4216714d, 32'hc0fb7bd0} /* (21, 0, 14) {real, imag} */,
  {32'hc13b46ba, 32'hc1d0075f} /* (21, 0, 13) {real, imag} */,
  {32'h423f9fc9, 32'h427f0f22} /* (21, 0, 12) {real, imag} */,
  {32'hc2144a57, 32'hc2722322} /* (21, 0, 11) {real, imag} */,
  {32'h417a010b, 32'h431d13b6} /* (21, 0, 10) {real, imag} */,
  {32'h4289386d, 32'h40a366ac} /* (21, 0, 9) {real, imag} */,
  {32'hc1c182df, 32'hbfee5680} /* (21, 0, 8) {real, imag} */,
  {32'hc1aa5fd4, 32'hc2af723a} /* (21, 0, 7) {real, imag} */,
  {32'hc2745329, 32'h41dc03bc} /* (21, 0, 6) {real, imag} */,
  {32'h42a63412, 32'h41e3c34c} /* (21, 0, 5) {real, imag} */,
  {32'hc18babf0, 32'h432716b9} /* (21, 0, 4) {real, imag} */,
  {32'h43619e64, 32'hc19b2a64} /* (21, 0, 3) {real, imag} */,
  {32'h4380d046, 32'h44430249} /* (21, 0, 2) {real, imag} */,
  {32'hc56c4589, 32'hc545a4e8} /* (21, 0, 1) {real, imag} */,
  {32'hc5aa0cf8, 32'h00000000} /* (21, 0, 0) {real, imag} */,
  {32'hc581f7a3, 32'h450f1b06} /* (20, 31, 31) {real, imag} */,
  {32'h4449e391, 32'hc40f5c30} /* (20, 31, 30) {real, imag} */,
  {32'h4291581d, 32'hc215fb03} /* (20, 31, 29) {real, imag} */,
  {32'hc291a406, 32'h4142bbc0} /* (20, 31, 28) {real, imag} */,
  {32'h42a225ba, 32'h41baf6c8} /* (20, 31, 27) {real, imag} */,
  {32'hc184ed28, 32'h4198626b} /* (20, 31, 26) {real, imag} */,
  {32'h40ed9738, 32'h42116b0a} /* (20, 31, 25) {real, imag} */,
  {32'h41957de6, 32'hc1bb7f6c} /* (20, 31, 24) {real, imag} */,
  {32'hbfa4f400, 32'hc2a12106} /* (20, 31, 23) {real, imag} */,
  {32'h42496a91, 32'h3e32ea00} /* (20, 31, 22) {real, imag} */,
  {32'hc1032df8, 32'h42909272} /* (20, 31, 21) {real, imag} */,
  {32'h4206063e, 32'h41b81177} /* (20, 31, 20) {real, imag} */,
  {32'hc15c13c4, 32'hc1b2fe69} /* (20, 31, 19) {real, imag} */,
  {32'h40a36522, 32'hc2150e8a} /* (20, 31, 18) {real, imag} */,
  {32'hc18ffed4, 32'hbfd03a00} /* (20, 31, 17) {real, imag} */,
  {32'h3ef47040, 32'h00000000} /* (20, 31, 16) {real, imag} */,
  {32'hc18ffed4, 32'h3fd03a00} /* (20, 31, 15) {real, imag} */,
  {32'h40a36522, 32'h42150e8a} /* (20, 31, 14) {real, imag} */,
  {32'hc15c13c4, 32'h41b2fe69} /* (20, 31, 13) {real, imag} */,
  {32'h4206063e, 32'hc1b81177} /* (20, 31, 12) {real, imag} */,
  {32'hc1032df8, 32'hc2909272} /* (20, 31, 11) {real, imag} */,
  {32'h42496a91, 32'hbe32ea00} /* (20, 31, 10) {real, imag} */,
  {32'hbfa4f400, 32'h42a12106} /* (20, 31, 9) {real, imag} */,
  {32'h41957de6, 32'h41bb7f6c} /* (20, 31, 8) {real, imag} */,
  {32'h40ed9738, 32'hc2116b0a} /* (20, 31, 7) {real, imag} */,
  {32'hc184ed28, 32'hc198626b} /* (20, 31, 6) {real, imag} */,
  {32'h42a225ba, 32'hc1baf6c8} /* (20, 31, 5) {real, imag} */,
  {32'hc291a406, 32'hc142bbc0} /* (20, 31, 4) {real, imag} */,
  {32'h4291581d, 32'h4215fb03} /* (20, 31, 3) {real, imag} */,
  {32'h4449e391, 32'h440f5c30} /* (20, 31, 2) {real, imag} */,
  {32'hc581f7a3, 32'hc50f1b06} /* (20, 31, 1) {real, imag} */,
  {32'hc5a31735, 32'h00000000} /* (20, 31, 0) {real, imag} */,
  {32'hc59923b2, 32'h44efb914} /* (20, 30, 31) {real, imag} */,
  {32'h44ab1562, 32'hc3e4ea26} /* (20, 30, 30) {real, imag} */,
  {32'h40707e90, 32'hc2202925} /* (20, 30, 29) {real, imag} */,
  {32'hc2200f71, 32'h43060458} /* (20, 30, 28) {real, imag} */,
  {32'h43326358, 32'h3f21cc70} /* (20, 30, 27) {real, imag} */,
  {32'hc1379acc, 32'hc215f178} /* (20, 30, 26) {real, imag} */,
  {32'hc0623a80, 32'h40294fd8} /* (20, 30, 25) {real, imag} */,
  {32'hc23b8f22, 32'hc154ed2a} /* (20, 30, 24) {real, imag} */,
  {32'hc2072a2c, 32'h4298ae31} /* (20, 30, 23) {real, imag} */,
  {32'h422d5c4f, 32'hc1314160} /* (20, 30, 22) {real, imag} */,
  {32'h424cea78, 32'hc145b672} /* (20, 30, 21) {real, imag} */,
  {32'h40e24e88, 32'hc219581a} /* (20, 30, 20) {real, imag} */,
  {32'hc2b5e9c8, 32'hc1db51d3} /* (20, 30, 19) {real, imag} */,
  {32'h42a87a94, 32'hc25f1b52} /* (20, 30, 18) {real, imag} */,
  {32'hc215b250, 32'h42540760} /* (20, 30, 17) {real, imag} */,
  {32'h427bd52e, 32'h00000000} /* (20, 30, 16) {real, imag} */,
  {32'hc215b250, 32'hc2540760} /* (20, 30, 15) {real, imag} */,
  {32'h42a87a94, 32'h425f1b52} /* (20, 30, 14) {real, imag} */,
  {32'hc2b5e9c8, 32'h41db51d3} /* (20, 30, 13) {real, imag} */,
  {32'h40e24e88, 32'h4219581a} /* (20, 30, 12) {real, imag} */,
  {32'h424cea78, 32'h4145b672} /* (20, 30, 11) {real, imag} */,
  {32'h422d5c4f, 32'h41314160} /* (20, 30, 10) {real, imag} */,
  {32'hc2072a2c, 32'hc298ae31} /* (20, 30, 9) {real, imag} */,
  {32'hc23b8f22, 32'h4154ed2a} /* (20, 30, 8) {real, imag} */,
  {32'hc0623a80, 32'hc0294fd8} /* (20, 30, 7) {real, imag} */,
  {32'hc1379acc, 32'h4215f178} /* (20, 30, 6) {real, imag} */,
  {32'h43326358, 32'hbf21cc70} /* (20, 30, 5) {real, imag} */,
  {32'hc2200f71, 32'hc3060458} /* (20, 30, 4) {real, imag} */,
  {32'h40707e90, 32'h42202925} /* (20, 30, 3) {real, imag} */,
  {32'h44ab1562, 32'h43e4ea26} /* (20, 30, 2) {real, imag} */,
  {32'hc59923b2, 32'hc4efb914} /* (20, 30, 1) {real, imag} */,
  {32'hc5a79342, 32'h00000000} /* (20, 30, 0) {real, imag} */,
  {32'hc59f4b31, 32'h44d4e3ea} /* (20, 29, 31) {real, imag} */,
  {32'h44bf427a, 32'hc3af812b} /* (20, 29, 30) {real, imag} */,
  {32'h420e71ed, 32'hc260ea7a} /* (20, 29, 29) {real, imag} */,
  {32'hc396abaa, 32'h42bb02e2} /* (20, 29, 28) {real, imag} */,
  {32'h42cea7ad, 32'hc24bd0af} /* (20, 29, 27) {real, imag} */,
  {32'hc1a5ec60, 32'hc22b4360} /* (20, 29, 26) {real, imag} */,
  {32'h41a4d43b, 32'h429b2905} /* (20, 29, 25) {real, imag} */,
  {32'h427293f4, 32'h4120e7d4} /* (20, 29, 24) {real, imag} */,
  {32'hc22640d5, 32'hc2825a2e} /* (20, 29, 23) {real, imag} */,
  {32'hc271a449, 32'h42be698c} /* (20, 29, 22) {real, imag} */,
  {32'h42029790, 32'hc2ad5b07} /* (20, 29, 21) {real, imag} */,
  {32'h4140c880, 32'hc23ca56e} /* (20, 29, 20) {real, imag} */,
  {32'h404cfeec, 32'h41de577c} /* (20, 29, 19) {real, imag} */,
  {32'h41321158, 32'h41384f70} /* (20, 29, 18) {real, imag} */,
  {32'h40d381c0, 32'hc1118934} /* (20, 29, 17) {real, imag} */,
  {32'hc2a849e8, 32'h00000000} /* (20, 29, 16) {real, imag} */,
  {32'h40d381c0, 32'h41118934} /* (20, 29, 15) {real, imag} */,
  {32'h41321158, 32'hc1384f70} /* (20, 29, 14) {real, imag} */,
  {32'h404cfeec, 32'hc1de577c} /* (20, 29, 13) {real, imag} */,
  {32'h4140c880, 32'h423ca56e} /* (20, 29, 12) {real, imag} */,
  {32'h42029790, 32'h42ad5b07} /* (20, 29, 11) {real, imag} */,
  {32'hc271a449, 32'hc2be698c} /* (20, 29, 10) {real, imag} */,
  {32'hc22640d5, 32'h42825a2e} /* (20, 29, 9) {real, imag} */,
  {32'h427293f4, 32'hc120e7d4} /* (20, 29, 8) {real, imag} */,
  {32'h41a4d43b, 32'hc29b2905} /* (20, 29, 7) {real, imag} */,
  {32'hc1a5ec60, 32'h422b4360} /* (20, 29, 6) {real, imag} */,
  {32'h42cea7ad, 32'h424bd0af} /* (20, 29, 5) {real, imag} */,
  {32'hc396abaa, 32'hc2bb02e2} /* (20, 29, 4) {real, imag} */,
  {32'h420e71ed, 32'h4260ea7a} /* (20, 29, 3) {real, imag} */,
  {32'h44bf427a, 32'h43af812b} /* (20, 29, 2) {real, imag} */,
  {32'hc59f4b31, 32'hc4d4e3ea} /* (20, 29, 1) {real, imag} */,
  {32'hc5a6bc94, 32'h00000000} /* (20, 29, 0) {real, imag} */,
  {32'hc5a3a2ea, 32'h44b5e290} /* (20, 28, 31) {real, imag} */,
  {32'h44de483e, 32'hc3fcf94b} /* (20, 28, 30) {real, imag} */,
  {32'h41c7de02, 32'hc2471878} /* (20, 28, 29) {real, imag} */,
  {32'hc3b3607f, 32'h42e1957f} /* (20, 28, 28) {real, imag} */,
  {32'h4299e8aa, 32'hc290c1e6} /* (20, 28, 27) {real, imag} */,
  {32'h42c93618, 32'hc21d05fb} /* (20, 28, 26) {real, imag} */,
  {32'hc30699b5, 32'h426e2428} /* (20, 28, 25) {real, imag} */,
  {32'hc245c037, 32'hc2dcdb7a} /* (20, 28, 24) {real, imag} */,
  {32'hc1f2690c, 32'hc23b7d0f} /* (20, 28, 23) {real, imag} */,
  {32'h411bf9c2, 32'hc183dd6a} /* (20, 28, 22) {real, imag} */,
  {32'h42c2f60d, 32'h4202298a} /* (20, 28, 21) {real, imag} */,
  {32'hc10ac2f1, 32'hc21f0e84} /* (20, 28, 20) {real, imag} */,
  {32'h4207051b, 32'hc1d70c3c} /* (20, 28, 19) {real, imag} */,
  {32'h409b72e8, 32'h3f0d20f0} /* (20, 28, 18) {real, imag} */,
  {32'hc1b3bf93, 32'hbfc189e0} /* (20, 28, 17) {real, imag} */,
  {32'hc287ca1d, 32'h00000000} /* (20, 28, 16) {real, imag} */,
  {32'hc1b3bf93, 32'h3fc189e0} /* (20, 28, 15) {real, imag} */,
  {32'h409b72e8, 32'hbf0d20f0} /* (20, 28, 14) {real, imag} */,
  {32'h4207051b, 32'h41d70c3c} /* (20, 28, 13) {real, imag} */,
  {32'hc10ac2f1, 32'h421f0e84} /* (20, 28, 12) {real, imag} */,
  {32'h42c2f60d, 32'hc202298a} /* (20, 28, 11) {real, imag} */,
  {32'h411bf9c2, 32'h4183dd6a} /* (20, 28, 10) {real, imag} */,
  {32'hc1f2690c, 32'h423b7d0f} /* (20, 28, 9) {real, imag} */,
  {32'hc245c037, 32'h42dcdb7a} /* (20, 28, 8) {real, imag} */,
  {32'hc30699b5, 32'hc26e2428} /* (20, 28, 7) {real, imag} */,
  {32'h42c93618, 32'h421d05fb} /* (20, 28, 6) {real, imag} */,
  {32'h4299e8aa, 32'h4290c1e6} /* (20, 28, 5) {real, imag} */,
  {32'hc3b3607f, 32'hc2e1957f} /* (20, 28, 4) {real, imag} */,
  {32'h41c7de02, 32'h42471878} /* (20, 28, 3) {real, imag} */,
  {32'h44de483e, 32'h43fcf94b} /* (20, 28, 2) {real, imag} */,
  {32'hc5a3a2ea, 32'hc4b5e290} /* (20, 28, 1) {real, imag} */,
  {32'hc5ab9dbe, 32'h00000000} /* (20, 28, 0) {real, imag} */,
  {32'hc5a6a3a9, 32'h448ee9a7} /* (20, 27, 31) {real, imag} */,
  {32'h44e47f0d, 32'hc4034d18} /* (20, 27, 30) {real, imag} */,
  {32'h4205dc80, 32'h424fe343} /* (20, 27, 29) {real, imag} */,
  {32'hc3464c3a, 32'h42dae1c7} /* (20, 27, 28) {real, imag} */,
  {32'h4352cc03, 32'hc262975f} /* (20, 27, 27) {real, imag} */,
  {32'h42c6ab37, 32'hc29c27b2} /* (20, 27, 26) {real, imag} */,
  {32'hc2eb9638, 32'hc2d2b0da} /* (20, 27, 25) {real, imag} */,
  {32'hc2127d0c, 32'hc225296a} /* (20, 27, 24) {real, imag} */,
  {32'h42c9fc74, 32'h42b3c946} /* (20, 27, 23) {real, imag} */,
  {32'h42c3fe4c, 32'h414caad4} /* (20, 27, 22) {real, imag} */,
  {32'hc14c27d4, 32'hc1bdadf4} /* (20, 27, 21) {real, imag} */,
  {32'h409e9908, 32'h4269cb3e} /* (20, 27, 20) {real, imag} */,
  {32'h422faee0, 32'h41309b9e} /* (20, 27, 19) {real, imag} */,
  {32'hc1cab958, 32'hc228c4be} /* (20, 27, 18) {real, imag} */,
  {32'hc011bfe0, 32'hc1a8417c} /* (20, 27, 17) {real, imag} */,
  {32'h415d43b0, 32'h00000000} /* (20, 27, 16) {real, imag} */,
  {32'hc011bfe0, 32'h41a8417c} /* (20, 27, 15) {real, imag} */,
  {32'hc1cab958, 32'h4228c4be} /* (20, 27, 14) {real, imag} */,
  {32'h422faee0, 32'hc1309b9e} /* (20, 27, 13) {real, imag} */,
  {32'h409e9908, 32'hc269cb3e} /* (20, 27, 12) {real, imag} */,
  {32'hc14c27d4, 32'h41bdadf4} /* (20, 27, 11) {real, imag} */,
  {32'h42c3fe4c, 32'hc14caad4} /* (20, 27, 10) {real, imag} */,
  {32'h42c9fc74, 32'hc2b3c946} /* (20, 27, 9) {real, imag} */,
  {32'hc2127d0c, 32'h4225296a} /* (20, 27, 8) {real, imag} */,
  {32'hc2eb9638, 32'h42d2b0da} /* (20, 27, 7) {real, imag} */,
  {32'h42c6ab37, 32'h429c27b2} /* (20, 27, 6) {real, imag} */,
  {32'h4352cc03, 32'h4262975f} /* (20, 27, 5) {real, imag} */,
  {32'hc3464c3a, 32'hc2dae1c7} /* (20, 27, 4) {real, imag} */,
  {32'h4205dc80, 32'hc24fe343} /* (20, 27, 3) {real, imag} */,
  {32'h44e47f0d, 32'h44034d18} /* (20, 27, 2) {real, imag} */,
  {32'hc5a6a3a9, 32'hc48ee9a7} /* (20, 27, 1) {real, imag} */,
  {32'hc5af427e, 32'h00000000} /* (20, 27, 0) {real, imag} */,
  {32'hc5a17475, 32'h447077c4} /* (20, 26, 31) {real, imag} */,
  {32'h44ec44b8, 32'hc3e82b13} /* (20, 26, 30) {real, imag} */,
  {32'hc26e5a28, 32'h42823503} /* (20, 26, 29) {real, imag} */,
  {32'hc39cbca2, 32'h4254fd2e} /* (20, 26, 28) {real, imag} */,
  {32'h43943d7c, 32'hc2ea9b62} /* (20, 26, 27) {real, imag} */,
  {32'hc10abc33, 32'hc30d7558} /* (20, 26, 26) {real, imag} */,
  {32'hc1fc14f0, 32'hc100900c} /* (20, 26, 25) {real, imag} */,
  {32'h4150cb70, 32'hc246ce72} /* (20, 26, 24) {real, imag} */,
  {32'hc1165e94, 32'h42882f52} /* (20, 26, 23) {real, imag} */,
  {32'hc2f18fc2, 32'hc203bc76} /* (20, 26, 22) {real, imag} */,
  {32'h42b3999c, 32'h41b96b9f} /* (20, 26, 21) {real, imag} */,
  {32'hc180c544, 32'h4214d950} /* (20, 26, 20) {real, imag} */,
  {32'h40608900, 32'hc22dbd82} /* (20, 26, 19) {real, imag} */,
  {32'hc1547d74, 32'hc284168a} /* (20, 26, 18) {real, imag} */,
  {32'hc1067543, 32'h41da5004} /* (20, 26, 17) {real, imag} */,
  {32'hc283a642, 32'h00000000} /* (20, 26, 16) {real, imag} */,
  {32'hc1067543, 32'hc1da5004} /* (20, 26, 15) {real, imag} */,
  {32'hc1547d74, 32'h4284168a} /* (20, 26, 14) {real, imag} */,
  {32'h40608900, 32'h422dbd82} /* (20, 26, 13) {real, imag} */,
  {32'hc180c544, 32'hc214d950} /* (20, 26, 12) {real, imag} */,
  {32'h42b3999c, 32'hc1b96b9f} /* (20, 26, 11) {real, imag} */,
  {32'hc2f18fc2, 32'h4203bc76} /* (20, 26, 10) {real, imag} */,
  {32'hc1165e94, 32'hc2882f52} /* (20, 26, 9) {real, imag} */,
  {32'h4150cb70, 32'h4246ce72} /* (20, 26, 8) {real, imag} */,
  {32'hc1fc14f0, 32'h4100900c} /* (20, 26, 7) {real, imag} */,
  {32'hc10abc33, 32'h430d7558} /* (20, 26, 6) {real, imag} */,
  {32'h43943d7c, 32'h42ea9b62} /* (20, 26, 5) {real, imag} */,
  {32'hc39cbca2, 32'hc254fd2e} /* (20, 26, 4) {real, imag} */,
  {32'hc26e5a28, 32'hc2823503} /* (20, 26, 3) {real, imag} */,
  {32'h44ec44b8, 32'h43e82b13} /* (20, 26, 2) {real, imag} */,
  {32'hc5a17475, 32'hc47077c4} /* (20, 26, 1) {real, imag} */,
  {32'hc5a42c09, 32'h00000000} /* (20, 26, 0) {real, imag} */,
  {32'hc59683fd, 32'h443514d5} /* (20, 25, 31) {real, imag} */,
  {32'h44e20683, 32'hc3ccb132} /* (20, 25, 30) {real, imag} */,
  {32'h413d6dd8, 32'h4329368e} /* (20, 25, 29) {real, imag} */,
  {32'hc3a8fa3c, 32'h4299f6d5} /* (20, 25, 28) {real, imag} */,
  {32'h4387eab4, 32'hc34f7cfd} /* (20, 25, 27) {real, imag} */,
  {32'hc2e4a6b2, 32'hc2d36286} /* (20, 25, 26) {real, imag} */,
  {32'h422c23a2, 32'h40f5d3b8} /* (20, 25, 25) {real, imag} */,
  {32'h42b35f24, 32'hc14c56e0} /* (20, 25, 24) {real, imag} */,
  {32'h418a7214, 32'h4181e39a} /* (20, 25, 23) {real, imag} */,
  {32'hc297be5b, 32'h42d33f00} /* (20, 25, 22) {real, imag} */,
  {32'h42e4257e, 32'h41fc35ff} /* (20, 25, 21) {real, imag} */,
  {32'h409367c4, 32'hc244fb36} /* (20, 25, 20) {real, imag} */,
  {32'hc23a6dc9, 32'h417d6580} /* (20, 25, 19) {real, imag} */,
  {32'h41c7977b, 32'hc1ed5ef2} /* (20, 25, 18) {real, imag} */,
  {32'hc250ce93, 32'h427a8924} /* (20, 25, 17) {real, imag} */,
  {32'h418febaa, 32'h00000000} /* (20, 25, 16) {real, imag} */,
  {32'hc250ce93, 32'hc27a8924} /* (20, 25, 15) {real, imag} */,
  {32'h41c7977b, 32'h41ed5ef2} /* (20, 25, 14) {real, imag} */,
  {32'hc23a6dc9, 32'hc17d6580} /* (20, 25, 13) {real, imag} */,
  {32'h409367c4, 32'h4244fb36} /* (20, 25, 12) {real, imag} */,
  {32'h42e4257e, 32'hc1fc35ff} /* (20, 25, 11) {real, imag} */,
  {32'hc297be5b, 32'hc2d33f00} /* (20, 25, 10) {real, imag} */,
  {32'h418a7214, 32'hc181e39a} /* (20, 25, 9) {real, imag} */,
  {32'h42b35f24, 32'h414c56e0} /* (20, 25, 8) {real, imag} */,
  {32'h422c23a2, 32'hc0f5d3b8} /* (20, 25, 7) {real, imag} */,
  {32'hc2e4a6b2, 32'h42d36286} /* (20, 25, 6) {real, imag} */,
  {32'h4387eab4, 32'h434f7cfd} /* (20, 25, 5) {real, imag} */,
  {32'hc3a8fa3c, 32'hc299f6d5} /* (20, 25, 4) {real, imag} */,
  {32'h413d6dd8, 32'hc329368e} /* (20, 25, 3) {real, imag} */,
  {32'h44e20683, 32'h43ccb132} /* (20, 25, 2) {real, imag} */,
  {32'hc59683fd, 32'hc43514d5} /* (20, 25, 1) {real, imag} */,
  {32'hc5970893, 32'h00000000} /* (20, 25, 0) {real, imag} */,
  {32'hc583e6e4, 32'h43c9f4bc} /* (20, 24, 31) {real, imag} */,
  {32'h44d38d6e, 32'hc3e5e0ef} /* (20, 24, 30) {real, imag} */,
  {32'hc266524e, 32'h40a399b8} /* (20, 24, 29) {real, imag} */,
  {32'hc3905998, 32'h41345bca} /* (20, 24, 28) {real, imag} */,
  {32'h43538bbd, 32'hc311bb7c} /* (20, 24, 27) {real, imag} */,
  {32'h4281d84c, 32'hc2c6651a} /* (20, 24, 26) {real, imag} */,
  {32'hc1a78d33, 32'h4252efb8} /* (20, 24, 25) {real, imag} */,
  {32'h429d11e3, 32'hc06c9380} /* (20, 24, 24) {real, imag} */,
  {32'h4203d01e, 32'h41c2af9a} /* (20, 24, 23) {real, imag} */,
  {32'hc1e32ff8, 32'h42d42942} /* (20, 24, 22) {real, imag} */,
  {32'hc262635c, 32'hc2636df3} /* (20, 24, 21) {real, imag} */,
  {32'hc310be86, 32'hc2895bf9} /* (20, 24, 20) {real, imag} */,
  {32'h4280979f, 32'hc28b7a39} /* (20, 24, 19) {real, imag} */,
  {32'hc03d8bb4, 32'h425951fe} /* (20, 24, 18) {real, imag} */,
  {32'hc2885d47, 32'h427f3145} /* (20, 24, 17) {real, imag} */,
  {32'hc213a6ec, 32'h00000000} /* (20, 24, 16) {real, imag} */,
  {32'hc2885d47, 32'hc27f3145} /* (20, 24, 15) {real, imag} */,
  {32'hc03d8bb4, 32'hc25951fe} /* (20, 24, 14) {real, imag} */,
  {32'h4280979f, 32'h428b7a39} /* (20, 24, 13) {real, imag} */,
  {32'hc310be86, 32'h42895bf9} /* (20, 24, 12) {real, imag} */,
  {32'hc262635c, 32'h42636df3} /* (20, 24, 11) {real, imag} */,
  {32'hc1e32ff8, 32'hc2d42942} /* (20, 24, 10) {real, imag} */,
  {32'h4203d01e, 32'hc1c2af9a} /* (20, 24, 9) {real, imag} */,
  {32'h429d11e3, 32'h406c9380} /* (20, 24, 8) {real, imag} */,
  {32'hc1a78d33, 32'hc252efb8} /* (20, 24, 7) {real, imag} */,
  {32'h4281d84c, 32'h42c6651a} /* (20, 24, 6) {real, imag} */,
  {32'h43538bbd, 32'h4311bb7c} /* (20, 24, 5) {real, imag} */,
  {32'hc3905998, 32'hc1345bca} /* (20, 24, 4) {real, imag} */,
  {32'hc266524e, 32'hc0a399b8} /* (20, 24, 3) {real, imag} */,
  {32'h44d38d6e, 32'h43e5e0ef} /* (20, 24, 2) {real, imag} */,
  {32'hc583e6e4, 32'hc3c9f4bc} /* (20, 24, 1) {real, imag} */,
  {32'hc5879053, 32'h00000000} /* (20, 24, 0) {real, imag} */,
  {32'hc5572b0a, 32'h439b6524} /* (20, 23, 31) {real, imag} */,
  {32'h44b478e9, 32'hc3ccb476} /* (20, 23, 30) {real, imag} */,
  {32'hc2bf1738, 32'hc2622f9c} /* (20, 23, 29) {real, imag} */,
  {32'hc369b93c, 32'hc202c8be} /* (20, 23, 28) {real, imag} */,
  {32'h4396b4e4, 32'hc3008958} /* (20, 23, 27) {real, imag} */,
  {32'hc29bc844, 32'hc2ab12b2} /* (20, 23, 26) {real, imag} */,
  {32'hc210dad0, 32'h40a0e860} /* (20, 23, 25) {real, imag} */,
  {32'h41b2443c, 32'hc2d4ad54} /* (20, 23, 24) {real, imag} */,
  {32'hc29712c1, 32'h42be1690} /* (20, 23, 23) {real, imag} */,
  {32'h42efc4d0, 32'hc1c0fccd} /* (20, 23, 22) {real, imag} */,
  {32'hc22c12a2, 32'hc2d35ef9} /* (20, 23, 21) {real, imag} */,
  {32'h4181480c, 32'h41961914} /* (20, 23, 20) {real, imag} */,
  {32'h4173dfab, 32'hc26f0d4c} /* (20, 23, 19) {real, imag} */,
  {32'h42137962, 32'hc20bcd9f} /* (20, 23, 18) {real, imag} */,
  {32'h41ccbdda, 32'h425a08d6} /* (20, 23, 17) {real, imag} */,
  {32'h41a60664, 32'h00000000} /* (20, 23, 16) {real, imag} */,
  {32'h41ccbdda, 32'hc25a08d6} /* (20, 23, 15) {real, imag} */,
  {32'h42137962, 32'h420bcd9f} /* (20, 23, 14) {real, imag} */,
  {32'h4173dfab, 32'h426f0d4c} /* (20, 23, 13) {real, imag} */,
  {32'h4181480c, 32'hc1961914} /* (20, 23, 12) {real, imag} */,
  {32'hc22c12a2, 32'h42d35ef9} /* (20, 23, 11) {real, imag} */,
  {32'h42efc4d0, 32'h41c0fccd} /* (20, 23, 10) {real, imag} */,
  {32'hc29712c1, 32'hc2be1690} /* (20, 23, 9) {real, imag} */,
  {32'h41b2443c, 32'h42d4ad54} /* (20, 23, 8) {real, imag} */,
  {32'hc210dad0, 32'hc0a0e860} /* (20, 23, 7) {real, imag} */,
  {32'hc29bc844, 32'h42ab12b2} /* (20, 23, 6) {real, imag} */,
  {32'h4396b4e4, 32'h43008958} /* (20, 23, 5) {real, imag} */,
  {32'hc369b93c, 32'h4202c8be} /* (20, 23, 4) {real, imag} */,
  {32'hc2bf1738, 32'h42622f9c} /* (20, 23, 3) {real, imag} */,
  {32'h44b478e9, 32'h43ccb476} /* (20, 23, 2) {real, imag} */,
  {32'hc5572b0a, 32'hc39b6524} /* (20, 23, 1) {real, imag} */,
  {32'hc55e9efb, 32'h00000000} /* (20, 23, 0) {real, imag} */,
  {32'hc51dcdbd, 32'h433bd170} /* (20, 22, 31) {real, imag} */,
  {32'h4480ea52, 32'hc39d36ad} /* (20, 22, 30) {real, imag} */,
  {32'hbf3f77c0, 32'h423ad6a0} /* (20, 22, 29) {real, imag} */,
  {32'hc39aebbb, 32'hc22c4468} /* (20, 22, 28) {real, imag} */,
  {32'h4392265a, 32'hc323cb96} /* (20, 22, 27) {real, imag} */,
  {32'hc23c32c0, 32'h4035f088} /* (20, 22, 26) {real, imag} */,
  {32'hc1641fec, 32'hc1b4b2a0} /* (20, 22, 25) {real, imag} */,
  {32'hc0a02d00, 32'hc2f06dd8} /* (20, 22, 24) {real, imag} */,
  {32'hc2828144, 32'h4232134b} /* (20, 22, 23) {real, imag} */,
  {32'hc0555f38, 32'hc20314fd} /* (20, 22, 22) {real, imag} */,
  {32'h40848fc0, 32'hc28fadd2} /* (20, 22, 21) {real, imag} */,
  {32'h427694d8, 32'hc1fcf21f} /* (20, 22, 20) {real, imag} */,
  {32'h41ff8fde, 32'hc1785a80} /* (20, 22, 19) {real, imag} */,
  {32'h41de4028, 32'hc0913560} /* (20, 22, 18) {real, imag} */,
  {32'h424297ce, 32'hc238be40} /* (20, 22, 17) {real, imag} */,
  {32'h429d4442, 32'h00000000} /* (20, 22, 16) {real, imag} */,
  {32'h424297ce, 32'h4238be40} /* (20, 22, 15) {real, imag} */,
  {32'h41de4028, 32'h40913560} /* (20, 22, 14) {real, imag} */,
  {32'h41ff8fde, 32'h41785a80} /* (20, 22, 13) {real, imag} */,
  {32'h427694d8, 32'h41fcf21f} /* (20, 22, 12) {real, imag} */,
  {32'h40848fc0, 32'h428fadd2} /* (20, 22, 11) {real, imag} */,
  {32'hc0555f38, 32'h420314fd} /* (20, 22, 10) {real, imag} */,
  {32'hc2828144, 32'hc232134b} /* (20, 22, 9) {real, imag} */,
  {32'hc0a02d00, 32'h42f06dd8} /* (20, 22, 8) {real, imag} */,
  {32'hc1641fec, 32'h41b4b2a0} /* (20, 22, 7) {real, imag} */,
  {32'hc23c32c0, 32'hc035f088} /* (20, 22, 6) {real, imag} */,
  {32'h4392265a, 32'h4323cb96} /* (20, 22, 5) {real, imag} */,
  {32'hc39aebbb, 32'h422c4468} /* (20, 22, 4) {real, imag} */,
  {32'hbf3f77c0, 32'hc23ad6a0} /* (20, 22, 3) {real, imag} */,
  {32'h4480ea52, 32'h439d36ad} /* (20, 22, 2) {real, imag} */,
  {32'hc51dcdbd, 32'hc33bd170} /* (20, 22, 1) {real, imag} */,
  {32'hc51d4479, 32'h00000000} /* (20, 22, 0) {real, imag} */,
  {32'hc46624a5, 32'h42792000} /* (20, 21, 31) {real, imag} */,
  {32'h43a303a8, 32'hc2df662e} /* (20, 21, 30) {real, imag} */,
  {32'hc29a3b10, 32'h434f760a} /* (20, 21, 29) {real, imag} */,
  {32'hc2ab100d, 32'hc2591a4e} /* (20, 21, 28) {real, imag} */,
  {32'h42e6b612, 32'h4166375c} /* (20, 21, 27) {real, imag} */,
  {32'h3f963878, 32'hbfa17130} /* (20, 21, 26) {real, imag} */,
  {32'h41ad6255, 32'hc296a914} /* (20, 21, 25) {real, imag} */,
  {32'hc190001c, 32'hc22d366c} /* (20, 21, 24) {real, imag} */,
  {32'h42967dc7, 32'h41aaee82} /* (20, 21, 23) {real, imag} */,
  {32'hc30cf9d2, 32'hc276edcb} /* (20, 21, 22) {real, imag} */,
  {32'h42a8563e, 32'hc2882df3} /* (20, 21, 21) {real, imag} */,
  {32'h43313ba6, 32'h4150a1c0} /* (20, 21, 20) {real, imag} */,
  {32'hc24e240e, 32'h412c9409} /* (20, 21, 19) {real, imag} */,
  {32'h4208be72, 32'h42c30613} /* (20, 21, 18) {real, imag} */,
  {32'hc1953eb3, 32'hc1f865b8} /* (20, 21, 17) {real, imag} */,
  {32'hc2e592c7, 32'h00000000} /* (20, 21, 16) {real, imag} */,
  {32'hc1953eb3, 32'h41f865b8} /* (20, 21, 15) {real, imag} */,
  {32'h4208be72, 32'hc2c30613} /* (20, 21, 14) {real, imag} */,
  {32'hc24e240e, 32'hc12c9409} /* (20, 21, 13) {real, imag} */,
  {32'h43313ba6, 32'hc150a1c0} /* (20, 21, 12) {real, imag} */,
  {32'h42a8563e, 32'h42882df3} /* (20, 21, 11) {real, imag} */,
  {32'hc30cf9d2, 32'h4276edcb} /* (20, 21, 10) {real, imag} */,
  {32'h42967dc7, 32'hc1aaee82} /* (20, 21, 9) {real, imag} */,
  {32'hc190001c, 32'h422d366c} /* (20, 21, 8) {real, imag} */,
  {32'h41ad6255, 32'h4296a914} /* (20, 21, 7) {real, imag} */,
  {32'h3f963878, 32'h3fa17130} /* (20, 21, 6) {real, imag} */,
  {32'h42e6b612, 32'hc166375c} /* (20, 21, 5) {real, imag} */,
  {32'hc2ab100d, 32'h42591a4e} /* (20, 21, 4) {real, imag} */,
  {32'hc29a3b10, 32'hc34f760a} /* (20, 21, 3) {real, imag} */,
  {32'h43a303a8, 32'h42df662e} /* (20, 21, 2) {real, imag} */,
  {32'hc46624a5, 32'hc2792000} /* (20, 21, 1) {real, imag} */,
  {32'hc49957e8, 32'h00000000} /* (20, 21, 0) {real, imag} */,
  {32'h44979ad2, 32'hc3a9ad46} /* (20, 20, 31) {real, imag} */,
  {32'hc3f5db26, 32'h42a5b4f0} /* (20, 20, 30) {real, imag} */,
  {32'hc22932aa, 32'h4215a9fe} /* (20, 20, 29) {real, imag} */,
  {32'h3fa942c0, 32'hc35300c4} /* (20, 20, 28) {real, imag} */,
  {32'hc2808ae4, 32'h42a02f62} /* (20, 20, 27) {real, imag} */,
  {32'h42665e61, 32'hc209d682} /* (20, 20, 26) {real, imag} */,
  {32'hc17f94ca, 32'hc2c2a7fd} /* (20, 20, 25) {real, imag} */,
  {32'hc34cf254, 32'h42e88649} /* (20, 20, 24) {real, imag} */,
  {32'hc2a16fa2, 32'hc22bb0bf} /* (20, 20, 23) {real, imag} */,
  {32'hc285f384, 32'hc2af42fc} /* (20, 20, 22) {real, imag} */,
  {32'h41db0fad, 32'h429a0ada} /* (20, 20, 21) {real, imag} */,
  {32'h41888282, 32'h41eaa86c} /* (20, 20, 20) {real, imag} */,
  {32'h4119f296, 32'h4199d7d6} /* (20, 20, 19) {real, imag} */,
  {32'h4185076e, 32'h4195b1ae} /* (20, 20, 18) {real, imag} */,
  {32'hc1a1091d, 32'hc0cb01f4} /* (20, 20, 17) {real, imag} */,
  {32'h4199fef7, 32'h00000000} /* (20, 20, 16) {real, imag} */,
  {32'hc1a1091d, 32'h40cb01f4} /* (20, 20, 15) {real, imag} */,
  {32'h4185076e, 32'hc195b1ae} /* (20, 20, 14) {real, imag} */,
  {32'h4119f296, 32'hc199d7d6} /* (20, 20, 13) {real, imag} */,
  {32'h41888282, 32'hc1eaa86c} /* (20, 20, 12) {real, imag} */,
  {32'h41db0fad, 32'hc29a0ada} /* (20, 20, 11) {real, imag} */,
  {32'hc285f384, 32'h42af42fc} /* (20, 20, 10) {real, imag} */,
  {32'hc2a16fa2, 32'h422bb0bf} /* (20, 20, 9) {real, imag} */,
  {32'hc34cf254, 32'hc2e88649} /* (20, 20, 8) {real, imag} */,
  {32'hc17f94ca, 32'h42c2a7fd} /* (20, 20, 7) {real, imag} */,
  {32'h42665e61, 32'h4209d682} /* (20, 20, 6) {real, imag} */,
  {32'hc2808ae4, 32'hc2a02f62} /* (20, 20, 5) {real, imag} */,
  {32'h3fa942c0, 32'h435300c4} /* (20, 20, 4) {real, imag} */,
  {32'hc22932aa, 32'hc215a9fe} /* (20, 20, 3) {real, imag} */,
  {32'hc3f5db26, 32'hc2a5b4f0} /* (20, 20, 2) {real, imag} */,
  {32'h44979ad2, 32'h43a9ad46} /* (20, 20, 1) {real, imag} */,
  {32'h43978e10, 32'h00000000} /* (20, 20, 0) {real, imag} */,
  {32'h4529951d, 32'hc40a6b8e} /* (20, 19, 31) {real, imag} */,
  {32'hc4858203, 32'h43181488} /* (20, 19, 30) {real, imag} */,
  {32'h4317ce9b, 32'h42ded765} /* (20, 19, 29) {real, imag} */,
  {32'h43070d9b, 32'hc29cc6d9} /* (20, 19, 28) {real, imag} */,
  {32'hc341a794, 32'h42816396} /* (20, 19, 27) {real, imag} */,
  {32'hc2689051, 32'h42aa467d} /* (20, 19, 26) {real, imag} */,
  {32'h42daa742, 32'h41b4d26a} /* (20, 19, 25) {real, imag} */,
  {32'h42056008, 32'h42df8f86} /* (20, 19, 24) {real, imag} */,
  {32'hc2a5aa88, 32'h41d7e176} /* (20, 19, 23) {real, imag} */,
  {32'h4246894d, 32'hc1282950} /* (20, 19, 22) {real, imag} */,
  {32'h4186d96e, 32'h4297c782} /* (20, 19, 21) {real, imag} */,
  {32'hc2caac53, 32'h4256c6ee} /* (20, 19, 20) {real, imag} */,
  {32'hc21aa3fe, 32'hc251ba43} /* (20, 19, 19) {real, imag} */,
  {32'h412d22f0, 32'h41edeec2} /* (20, 19, 18) {real, imag} */,
  {32'hc208be3d, 32'hc221f0ee} /* (20, 19, 17) {real, imag} */,
  {32'hc155914c, 32'h00000000} /* (20, 19, 16) {real, imag} */,
  {32'hc208be3d, 32'h4221f0ee} /* (20, 19, 15) {real, imag} */,
  {32'h412d22f0, 32'hc1edeec2} /* (20, 19, 14) {real, imag} */,
  {32'hc21aa3fe, 32'h4251ba43} /* (20, 19, 13) {real, imag} */,
  {32'hc2caac53, 32'hc256c6ee} /* (20, 19, 12) {real, imag} */,
  {32'h4186d96e, 32'hc297c782} /* (20, 19, 11) {real, imag} */,
  {32'h4246894d, 32'h41282950} /* (20, 19, 10) {real, imag} */,
  {32'hc2a5aa88, 32'hc1d7e176} /* (20, 19, 9) {real, imag} */,
  {32'h42056008, 32'hc2df8f86} /* (20, 19, 8) {real, imag} */,
  {32'h42daa742, 32'hc1b4d26a} /* (20, 19, 7) {real, imag} */,
  {32'hc2689051, 32'hc2aa467d} /* (20, 19, 6) {real, imag} */,
  {32'hc341a794, 32'hc2816396} /* (20, 19, 5) {real, imag} */,
  {32'h43070d9b, 32'h429cc6d9} /* (20, 19, 4) {real, imag} */,
  {32'h4317ce9b, 32'hc2ded765} /* (20, 19, 3) {real, imag} */,
  {32'hc4858203, 32'hc3181488} /* (20, 19, 2) {real, imag} */,
  {32'h4529951d, 32'h440a6b8e} /* (20, 19, 1) {real, imag} */,
  {32'h44a8feb5, 32'h00000000} /* (20, 19, 0) {real, imag} */,
  {32'h45651d40, 32'hc3f68438} /* (20, 18, 31) {real, imag} */,
  {32'hc4adab4c, 32'h438cf7ea} /* (20, 18, 30) {real, imag} */,
  {32'h4353a886, 32'h431d8a13} /* (20, 18, 29) {real, imag} */,
  {32'h42a7fea6, 32'hc2dc6c93} /* (20, 18, 28) {real, imag} */,
  {32'hc2f59b36, 32'h42dccec5} /* (20, 18, 27) {real, imag} */,
  {32'h41a061a8, 32'h41e8b7fe} /* (20, 18, 26) {real, imag} */,
  {32'h432d3066, 32'h42a2ca2f} /* (20, 18, 25) {real, imag} */,
  {32'h4235d6b5, 32'h4306027f} /* (20, 18, 24) {real, imag} */,
  {32'h425b0be7, 32'h41ad76c1} /* (20, 18, 23) {real, imag} */,
  {32'hc23e0081, 32'h42c8fda4} /* (20, 18, 22) {real, imag} */,
  {32'h42848772, 32'h42cf4a86} /* (20, 18, 21) {real, imag} */,
  {32'h431b7e11, 32'hc2a97d19} /* (20, 18, 20) {real, imag} */,
  {32'h4237010c, 32'h429b7400} /* (20, 18, 19) {real, imag} */,
  {32'h419b1f78, 32'h42a695c7} /* (20, 18, 18) {real, imag} */,
  {32'h4284f7b2, 32'hc2644420} /* (20, 18, 17) {real, imag} */,
  {32'hc0bf8818, 32'h00000000} /* (20, 18, 16) {real, imag} */,
  {32'h4284f7b2, 32'h42644420} /* (20, 18, 15) {real, imag} */,
  {32'h419b1f78, 32'hc2a695c7} /* (20, 18, 14) {real, imag} */,
  {32'h4237010c, 32'hc29b7400} /* (20, 18, 13) {real, imag} */,
  {32'h431b7e11, 32'h42a97d19} /* (20, 18, 12) {real, imag} */,
  {32'h42848772, 32'hc2cf4a86} /* (20, 18, 11) {real, imag} */,
  {32'hc23e0081, 32'hc2c8fda4} /* (20, 18, 10) {real, imag} */,
  {32'h425b0be7, 32'hc1ad76c1} /* (20, 18, 9) {real, imag} */,
  {32'h4235d6b5, 32'hc306027f} /* (20, 18, 8) {real, imag} */,
  {32'h432d3066, 32'hc2a2ca2f} /* (20, 18, 7) {real, imag} */,
  {32'h41a061a8, 32'hc1e8b7fe} /* (20, 18, 6) {real, imag} */,
  {32'hc2f59b36, 32'hc2dccec5} /* (20, 18, 5) {real, imag} */,
  {32'h42a7fea6, 32'h42dc6c93} /* (20, 18, 4) {real, imag} */,
  {32'h4353a886, 32'hc31d8a13} /* (20, 18, 3) {real, imag} */,
  {32'hc4adab4c, 32'hc38cf7ea} /* (20, 18, 2) {real, imag} */,
  {32'h45651d40, 32'h43f68438} /* (20, 18, 1) {real, imag} */,
  {32'h45136f46, 32'h00000000} /* (20, 18, 0) {real, imag} */,
  {32'h45853c97, 32'hc3e2edb0} /* (20, 17, 31) {real, imag} */,
  {32'hc4bd7904, 32'h4396b539} /* (20, 17, 30) {real, imag} */,
  {32'h417b6800, 32'h43348b58} /* (20, 17, 29) {real, imag} */,
  {32'h42f3b150, 32'h4119faa0} /* (20, 17, 28) {real, imag} */,
  {32'hc283637a, 32'h42c5c54d} /* (20, 17, 27) {real, imag} */,
  {32'hc20d0387, 32'h4257cb0c} /* (20, 17, 26) {real, imag} */,
  {32'h42b4d180, 32'hc25abf86} /* (20, 17, 25) {real, imag} */,
  {32'h41515d50, 32'h434bb49a} /* (20, 17, 24) {real, imag} */,
  {32'hc2572ce5, 32'h41c3d910} /* (20, 17, 23) {real, imag} */,
  {32'hc28884ae, 32'h42aec4df} /* (20, 17, 22) {real, imag} */,
  {32'hc19f473c, 32'hc1aa34fc} /* (20, 17, 21) {real, imag} */,
  {32'hc2f32930, 32'h420458fa} /* (20, 17, 20) {real, imag} */,
  {32'hc12b4166, 32'hc2091804} /* (20, 17, 19) {real, imag} */,
  {32'hc2d589d4, 32'h41944ae6} /* (20, 17, 18) {real, imag} */,
  {32'h41630888, 32'h42697dfd} /* (20, 17, 17) {real, imag} */,
  {32'hc13c6cd6, 32'h00000000} /* (20, 17, 16) {real, imag} */,
  {32'h41630888, 32'hc2697dfd} /* (20, 17, 15) {real, imag} */,
  {32'hc2d589d4, 32'hc1944ae6} /* (20, 17, 14) {real, imag} */,
  {32'hc12b4166, 32'h42091804} /* (20, 17, 13) {real, imag} */,
  {32'hc2f32930, 32'hc20458fa} /* (20, 17, 12) {real, imag} */,
  {32'hc19f473c, 32'h41aa34fc} /* (20, 17, 11) {real, imag} */,
  {32'hc28884ae, 32'hc2aec4df} /* (20, 17, 10) {real, imag} */,
  {32'hc2572ce5, 32'hc1c3d910} /* (20, 17, 9) {real, imag} */,
  {32'h41515d50, 32'hc34bb49a} /* (20, 17, 8) {real, imag} */,
  {32'h42b4d180, 32'h425abf86} /* (20, 17, 7) {real, imag} */,
  {32'hc20d0387, 32'hc257cb0c} /* (20, 17, 6) {real, imag} */,
  {32'hc283637a, 32'hc2c5c54d} /* (20, 17, 5) {real, imag} */,
  {32'h42f3b150, 32'hc119faa0} /* (20, 17, 4) {real, imag} */,
  {32'h417b6800, 32'hc3348b58} /* (20, 17, 3) {real, imag} */,
  {32'hc4bd7904, 32'hc396b539} /* (20, 17, 2) {real, imag} */,
  {32'h45853c97, 32'h43e2edb0} /* (20, 17, 1) {real, imag} */,
  {32'h45376323, 32'h00000000} /* (20, 17, 0) {real, imag} */,
  {32'h458c7d09, 32'hc3d91a60} /* (20, 16, 31) {real, imag} */,
  {32'hc4c4cc8f, 32'h43918204} /* (20, 16, 30) {real, imag} */,
  {32'hc2d577a0, 32'h4278213f} /* (20, 16, 29) {real, imag} */,
  {32'h437ce630, 32'h40f58c80} /* (20, 16, 28) {real, imag} */,
  {32'hc3333520, 32'h42d6b5be} /* (20, 16, 27) {real, imag} */,
  {32'hc27f2f84, 32'hc2b3b473} /* (20, 16, 26) {real, imag} */,
  {32'h42ee110f, 32'hc103017c} /* (20, 16, 25) {real, imag} */,
  {32'h40c92e6c, 32'h422d16b9} /* (20, 16, 24) {real, imag} */,
  {32'hc1942a8e, 32'h4109ed88} /* (20, 16, 23) {real, imag} */,
  {32'hc1fe20e9, 32'hc2b634a6} /* (20, 16, 22) {real, imag} */,
  {32'h413eae0e, 32'h41b1f20f} /* (20, 16, 21) {real, imag} */,
  {32'h418804ae, 32'h411c5570} /* (20, 16, 20) {real, imag} */,
  {32'h42a4f4c1, 32'h4217759f} /* (20, 16, 19) {real, imag} */,
  {32'hc05c1ca0, 32'hc12255b9} /* (20, 16, 18) {real, imag} */,
  {32'h4221fcb2, 32'hc21c8789} /* (20, 16, 17) {real, imag} */,
  {32'h402b3254, 32'h00000000} /* (20, 16, 16) {real, imag} */,
  {32'h4221fcb2, 32'h421c8789} /* (20, 16, 15) {real, imag} */,
  {32'hc05c1ca0, 32'h412255b9} /* (20, 16, 14) {real, imag} */,
  {32'h42a4f4c1, 32'hc217759f} /* (20, 16, 13) {real, imag} */,
  {32'h418804ae, 32'hc11c5570} /* (20, 16, 12) {real, imag} */,
  {32'h413eae0e, 32'hc1b1f20f} /* (20, 16, 11) {real, imag} */,
  {32'hc1fe20e9, 32'h42b634a6} /* (20, 16, 10) {real, imag} */,
  {32'hc1942a8e, 32'hc109ed88} /* (20, 16, 9) {real, imag} */,
  {32'h40c92e6c, 32'hc22d16b9} /* (20, 16, 8) {real, imag} */,
  {32'h42ee110f, 32'h4103017c} /* (20, 16, 7) {real, imag} */,
  {32'hc27f2f84, 32'h42b3b473} /* (20, 16, 6) {real, imag} */,
  {32'hc3333520, 32'hc2d6b5be} /* (20, 16, 5) {real, imag} */,
  {32'h437ce630, 32'hc0f58c80} /* (20, 16, 4) {real, imag} */,
  {32'hc2d577a0, 32'hc278213f} /* (20, 16, 3) {real, imag} */,
  {32'hc4c4cc8f, 32'hc3918204} /* (20, 16, 2) {real, imag} */,
  {32'h458c7d09, 32'h43d91a60} /* (20, 16, 1) {real, imag} */,
  {32'h454444fc, 32'h00000000} /* (20, 16, 0) {real, imag} */,
  {32'h458e8351, 32'hc3ce2fc8} /* (20, 15, 31) {real, imag} */,
  {32'hc4bcd816, 32'h43d1d735} /* (20, 15, 30) {real, imag} */,
  {32'hc2f2803c, 32'h419bc054} /* (20, 15, 29) {real, imag} */,
  {32'h4327e880, 32'hc32b6ff4} /* (20, 15, 28) {real, imag} */,
  {32'hc3a243a4, 32'h42dcd343} /* (20, 15, 27) {real, imag} */,
  {32'hc2b1d3c8, 32'hc2df68a8} /* (20, 15, 26) {real, imag} */,
  {32'hc2528f45, 32'hc2f60e25} /* (20, 15, 25) {real, imag} */,
  {32'hc324bf60, 32'h42c45794} /* (20, 15, 24) {real, imag} */,
  {32'h426b5afb, 32'hc29254f1} /* (20, 15, 23) {real, imag} */,
  {32'hc25aa450, 32'hc23293ca} /* (20, 15, 22) {real, imag} */,
  {32'h4293076a, 32'h419febb6} /* (20, 15, 21) {real, imag} */,
  {32'h4220e8d0, 32'hc2ace051} /* (20, 15, 20) {real, imag} */,
  {32'h411a2496, 32'hc1bd3ec8} /* (20, 15, 19) {real, imag} */,
  {32'h42222bd9, 32'h41bf5ee2} /* (20, 15, 18) {real, imag} */,
  {32'hc2d2cb81, 32'h425b949d} /* (20, 15, 17) {real, imag} */,
  {32'h3fa3c5a0, 32'h00000000} /* (20, 15, 16) {real, imag} */,
  {32'hc2d2cb81, 32'hc25b949d} /* (20, 15, 15) {real, imag} */,
  {32'h42222bd9, 32'hc1bf5ee2} /* (20, 15, 14) {real, imag} */,
  {32'h411a2496, 32'h41bd3ec8} /* (20, 15, 13) {real, imag} */,
  {32'h4220e8d0, 32'h42ace051} /* (20, 15, 12) {real, imag} */,
  {32'h4293076a, 32'hc19febb6} /* (20, 15, 11) {real, imag} */,
  {32'hc25aa450, 32'h423293ca} /* (20, 15, 10) {real, imag} */,
  {32'h426b5afb, 32'h429254f1} /* (20, 15, 9) {real, imag} */,
  {32'hc324bf60, 32'hc2c45794} /* (20, 15, 8) {real, imag} */,
  {32'hc2528f45, 32'h42f60e25} /* (20, 15, 7) {real, imag} */,
  {32'hc2b1d3c8, 32'h42df68a8} /* (20, 15, 6) {real, imag} */,
  {32'hc3a243a4, 32'hc2dcd343} /* (20, 15, 5) {real, imag} */,
  {32'h4327e880, 32'h432b6ff4} /* (20, 15, 4) {real, imag} */,
  {32'hc2f2803c, 32'hc19bc054} /* (20, 15, 3) {real, imag} */,
  {32'hc4bcd816, 32'hc3d1d735} /* (20, 15, 2) {real, imag} */,
  {32'h458e8351, 32'h43ce2fc8} /* (20, 15, 1) {real, imag} */,
  {32'h45411a7f, 32'h00000000} /* (20, 15, 0) {real, imag} */,
  {32'h45792a38, 32'hc3a14308} /* (20, 14, 31) {real, imag} */,
  {32'hc4c9684c, 32'h43a36ec6} /* (20, 14, 30) {real, imag} */,
  {32'hc1f37a40, 32'hc2b825ee} /* (20, 14, 29) {real, imag} */,
  {32'h43919f18, 32'hc2bb3cbb} /* (20, 14, 28) {real, imag} */,
  {32'hc361779f, 32'h42ffd84f} /* (20, 14, 27) {real, imag} */,
  {32'hc1e3b2e8, 32'h429937cc} /* (20, 14, 26) {real, imag} */,
  {32'h4201bec6, 32'hc23aa84e} /* (20, 14, 25) {real, imag} */,
  {32'hc29069c0, 32'h42bb8717} /* (20, 14, 24) {real, imag} */,
  {32'h420a23cd, 32'h41b8c603} /* (20, 14, 23) {real, imag} */,
  {32'hc21b9069, 32'hc1ea1210} /* (20, 14, 22) {real, imag} */,
  {32'hc286675e, 32'h412675ac} /* (20, 14, 21) {real, imag} */,
  {32'h42159a85, 32'hc0b878d0} /* (20, 14, 20) {real, imag} */,
  {32'hc304c135, 32'h41b061e9} /* (20, 14, 19) {real, imag} */,
  {32'hc2098c61, 32'h4211e26e} /* (20, 14, 18) {real, imag} */,
  {32'h41ad693a, 32'h41684c48} /* (20, 14, 17) {real, imag} */,
  {32'hc2426a76, 32'h00000000} /* (20, 14, 16) {real, imag} */,
  {32'h41ad693a, 32'hc1684c48} /* (20, 14, 15) {real, imag} */,
  {32'hc2098c61, 32'hc211e26e} /* (20, 14, 14) {real, imag} */,
  {32'hc304c135, 32'hc1b061e9} /* (20, 14, 13) {real, imag} */,
  {32'h42159a85, 32'h40b878d0} /* (20, 14, 12) {real, imag} */,
  {32'hc286675e, 32'hc12675ac} /* (20, 14, 11) {real, imag} */,
  {32'hc21b9069, 32'h41ea1210} /* (20, 14, 10) {real, imag} */,
  {32'h420a23cd, 32'hc1b8c603} /* (20, 14, 9) {real, imag} */,
  {32'hc29069c0, 32'hc2bb8717} /* (20, 14, 8) {real, imag} */,
  {32'h4201bec6, 32'h423aa84e} /* (20, 14, 7) {real, imag} */,
  {32'hc1e3b2e8, 32'hc29937cc} /* (20, 14, 6) {real, imag} */,
  {32'hc361779f, 32'hc2ffd84f} /* (20, 14, 5) {real, imag} */,
  {32'h43919f18, 32'h42bb3cbb} /* (20, 14, 4) {real, imag} */,
  {32'hc1f37a40, 32'h42b825ee} /* (20, 14, 3) {real, imag} */,
  {32'hc4c9684c, 32'hc3a36ec6} /* (20, 14, 2) {real, imag} */,
  {32'h45792a38, 32'h43a14308} /* (20, 14, 1) {real, imag} */,
  {32'h45334992, 32'h00000000} /* (20, 14, 0) {real, imag} */,
  {32'h454fb1af, 32'hc33fb158} /* (20, 13, 31) {real, imag} */,
  {32'hc4b3e6c1, 32'h43a8d8fa} /* (20, 13, 30) {real, imag} */,
  {32'hc1cb8412, 32'hc32cd8a2} /* (20, 13, 29) {real, imag} */,
  {32'h4380063a, 32'hc1b8d43c} /* (20, 13, 28) {real, imag} */,
  {32'hc38306dd, 32'h43400d53} /* (20, 13, 27) {real, imag} */,
  {32'h424c3225, 32'h41f21c6b} /* (20, 13, 26) {real, imag} */,
  {32'h4300dc35, 32'hc190dd66} /* (20, 13, 25) {real, imag} */,
  {32'h40dc05f4, 32'h41d4e8c8} /* (20, 13, 24) {real, imag} */,
  {32'hc2092fdf, 32'h42f08a3a} /* (20, 13, 23) {real, imag} */,
  {32'hc29f4419, 32'hc0d9cbd0} /* (20, 13, 22) {real, imag} */,
  {32'h423a1c83, 32'h429c66ac} /* (20, 13, 21) {real, imag} */,
  {32'h4243d776, 32'hc1b2de29} /* (20, 13, 20) {real, imag} */,
  {32'hc22288f8, 32'hc0215050} /* (20, 13, 19) {real, imag} */,
  {32'hc1b3f61e, 32'hc233c3d3} /* (20, 13, 18) {real, imag} */,
  {32'h40d7bc88, 32'hc1261ce8} /* (20, 13, 17) {real, imag} */,
  {32'h41f025c6, 32'h00000000} /* (20, 13, 16) {real, imag} */,
  {32'h40d7bc88, 32'h41261ce8} /* (20, 13, 15) {real, imag} */,
  {32'hc1b3f61e, 32'h4233c3d3} /* (20, 13, 14) {real, imag} */,
  {32'hc22288f8, 32'h40215050} /* (20, 13, 13) {real, imag} */,
  {32'h4243d776, 32'h41b2de29} /* (20, 13, 12) {real, imag} */,
  {32'h423a1c83, 32'hc29c66ac} /* (20, 13, 11) {real, imag} */,
  {32'hc29f4419, 32'h40d9cbd0} /* (20, 13, 10) {real, imag} */,
  {32'hc2092fdf, 32'hc2f08a3a} /* (20, 13, 9) {real, imag} */,
  {32'h40dc05f4, 32'hc1d4e8c8} /* (20, 13, 8) {real, imag} */,
  {32'h4300dc35, 32'h4190dd66} /* (20, 13, 7) {real, imag} */,
  {32'h424c3225, 32'hc1f21c6b} /* (20, 13, 6) {real, imag} */,
  {32'hc38306dd, 32'hc3400d53} /* (20, 13, 5) {real, imag} */,
  {32'h4380063a, 32'h41b8d43c} /* (20, 13, 4) {real, imag} */,
  {32'hc1cb8412, 32'h432cd8a2} /* (20, 13, 3) {real, imag} */,
  {32'hc4b3e6c1, 32'hc3a8d8fa} /* (20, 13, 2) {real, imag} */,
  {32'h454fb1af, 32'h433fb158} /* (20, 13, 1) {real, imag} */,
  {32'h451b4b16, 32'h00000000} /* (20, 13, 0) {real, imag} */,
  {32'h45134f91, 32'h431c064c} /* (20, 12, 31) {real, imag} */,
  {32'hc48f613c, 32'h439a0cce} /* (20, 12, 30) {real, imag} */,
  {32'h42f8eb0f, 32'hc33c99f2} /* (20, 12, 29) {real, imag} */,
  {32'h433183e8, 32'h420fc892} /* (20, 12, 28) {real, imag} */,
  {32'hc39dc1fc, 32'h42ec828e} /* (20, 12, 27) {real, imag} */,
  {32'h42997804, 32'h3f0039e0} /* (20, 12, 26) {real, imag} */,
  {32'hc2600d12, 32'hc347baee} /* (20, 12, 25) {real, imag} */,
  {32'hc1b4fd3c, 32'hc202fb1a} /* (20, 12, 24) {real, imag} */,
  {32'hc00bcfa0, 32'h427d9a35} /* (20, 12, 23) {real, imag} */,
  {32'hc21cce08, 32'hc0e9b868} /* (20, 12, 22) {real, imag} */,
  {32'h40005728, 32'h4291e484} /* (20, 12, 21) {real, imag} */,
  {32'hc2915ab4, 32'h41552e67} /* (20, 12, 20) {real, imag} */,
  {32'hc00bf176, 32'hc2719237} /* (20, 12, 19) {real, imag} */,
  {32'h4215ddaf, 32'h4287551a} /* (20, 12, 18) {real, imag} */,
  {32'hc1905f8d, 32'hc1a84e4f} /* (20, 12, 17) {real, imag} */,
  {32'h41341622, 32'h00000000} /* (20, 12, 16) {real, imag} */,
  {32'hc1905f8d, 32'h41a84e4f} /* (20, 12, 15) {real, imag} */,
  {32'h4215ddaf, 32'hc287551a} /* (20, 12, 14) {real, imag} */,
  {32'hc00bf176, 32'h42719237} /* (20, 12, 13) {real, imag} */,
  {32'hc2915ab4, 32'hc1552e67} /* (20, 12, 12) {real, imag} */,
  {32'h40005728, 32'hc291e484} /* (20, 12, 11) {real, imag} */,
  {32'hc21cce08, 32'h40e9b868} /* (20, 12, 10) {real, imag} */,
  {32'hc00bcfa0, 32'hc27d9a35} /* (20, 12, 9) {real, imag} */,
  {32'hc1b4fd3c, 32'h4202fb1a} /* (20, 12, 8) {real, imag} */,
  {32'hc2600d12, 32'h4347baee} /* (20, 12, 7) {real, imag} */,
  {32'h42997804, 32'hbf0039e0} /* (20, 12, 6) {real, imag} */,
  {32'hc39dc1fc, 32'hc2ec828e} /* (20, 12, 5) {real, imag} */,
  {32'h433183e8, 32'hc20fc892} /* (20, 12, 4) {real, imag} */,
  {32'h42f8eb0f, 32'h433c99f2} /* (20, 12, 3) {real, imag} */,
  {32'hc48f613c, 32'hc39a0cce} /* (20, 12, 2) {real, imag} */,
  {32'h45134f91, 32'hc31c064c} /* (20, 12, 1) {real, imag} */,
  {32'h44d59810, 32'h00000000} /* (20, 12, 0) {real, imag} */,
  {32'h44835a4e, 32'h43cc9598} /* (20, 11, 31) {real, imag} */,
  {32'hc4294aec, 32'hc2b88f8a} /* (20, 11, 30) {real, imag} */,
  {32'h419ab0c3, 32'hc2a56c40} /* (20, 11, 29) {real, imag} */,
  {32'h4303e8ea, 32'hc22c7606} /* (20, 11, 28) {real, imag} */,
  {32'hc357e4d3, 32'h430d2ca5} /* (20, 11, 27) {real, imag} */,
  {32'hc1cb92d0, 32'h422d02b2} /* (20, 11, 26) {real, imag} */,
  {32'h425d7328, 32'h4102eebc} /* (20, 11, 25) {real, imag} */,
  {32'hc3043dd0, 32'hc2a1e5f2} /* (20, 11, 24) {real, imag} */,
  {32'hc2e4f9dd, 32'hc28d1164} /* (20, 11, 23) {real, imag} */,
  {32'h41d1ff84, 32'h41a834d6} /* (20, 11, 22) {real, imag} */,
  {32'hc217f68f, 32'h41ce772d} /* (20, 11, 21) {real, imag} */,
  {32'h4297f033, 32'h422c6a47} /* (20, 11, 20) {real, imag} */,
  {32'hc23ff89a, 32'h41f7a73c} /* (20, 11, 19) {real, imag} */,
  {32'hc112df64, 32'h3f9ebb40} /* (20, 11, 18) {real, imag} */,
  {32'h420bf9b4, 32'h40ac057a} /* (20, 11, 17) {real, imag} */,
  {32'hc1190dc8, 32'h00000000} /* (20, 11, 16) {real, imag} */,
  {32'h420bf9b4, 32'hc0ac057a} /* (20, 11, 15) {real, imag} */,
  {32'hc112df64, 32'hbf9ebb40} /* (20, 11, 14) {real, imag} */,
  {32'hc23ff89a, 32'hc1f7a73c} /* (20, 11, 13) {real, imag} */,
  {32'h4297f033, 32'hc22c6a47} /* (20, 11, 12) {real, imag} */,
  {32'hc217f68f, 32'hc1ce772d} /* (20, 11, 11) {real, imag} */,
  {32'h41d1ff84, 32'hc1a834d6} /* (20, 11, 10) {real, imag} */,
  {32'hc2e4f9dd, 32'h428d1164} /* (20, 11, 9) {real, imag} */,
  {32'hc3043dd0, 32'h42a1e5f2} /* (20, 11, 8) {real, imag} */,
  {32'h425d7328, 32'hc102eebc} /* (20, 11, 7) {real, imag} */,
  {32'hc1cb92d0, 32'hc22d02b2} /* (20, 11, 6) {real, imag} */,
  {32'hc357e4d3, 32'hc30d2ca5} /* (20, 11, 5) {real, imag} */,
  {32'h4303e8ea, 32'h422c7606} /* (20, 11, 4) {real, imag} */,
  {32'h419ab0c3, 32'h42a56c40} /* (20, 11, 3) {real, imag} */,
  {32'hc4294aec, 32'h42b88f8a} /* (20, 11, 2) {real, imag} */,
  {32'h44835a4e, 32'hc3cc9598} /* (20, 11, 1) {real, imag} */,
  {32'h44401980, 32'h00000000} /* (20, 11, 0) {real, imag} */,
  {32'hc450a6b0, 32'h442fe9bc} /* (20, 10, 31) {real, imag} */,
  {32'h435d4704, 32'hc3644b56} /* (20, 10, 30) {real, imag} */,
  {32'hc1ca43ee, 32'hc2da1272} /* (20, 10, 29) {real, imag} */,
  {32'h42e60bcb, 32'hc23d6c0c} /* (20, 10, 28) {real, imag} */,
  {32'h413c4280, 32'hc215abc0} /* (20, 10, 27) {real, imag} */,
  {32'h41ff8bcc, 32'hc254fb56} /* (20, 10, 26) {real, imag} */,
  {32'hc1cd4bc0, 32'h42c0aaf4} /* (20, 10, 25) {real, imag} */,
  {32'h42d08b1c, 32'hc2257c50} /* (20, 10, 24) {real, imag} */,
  {32'h42baee3c, 32'hc0967da8} /* (20, 10, 23) {real, imag} */,
  {32'h42390a8c, 32'h42a01aaa} /* (20, 10, 22) {real, imag} */,
  {32'hc2d4a402, 32'h42ada9ee} /* (20, 10, 21) {real, imag} */,
  {32'hc07dcb20, 32'hc28a53fc} /* (20, 10, 20) {real, imag} */,
  {32'hc18b1dde, 32'h42772c26} /* (20, 10, 19) {real, imag} */,
  {32'hc0e0669a, 32'h420a6832} /* (20, 10, 18) {real, imag} */,
  {32'hc245515a, 32'hc0ba87c0} /* (20, 10, 17) {real, imag} */,
  {32'hc284d1a8, 32'h00000000} /* (20, 10, 16) {real, imag} */,
  {32'hc245515a, 32'h40ba87c0} /* (20, 10, 15) {real, imag} */,
  {32'hc0e0669a, 32'hc20a6832} /* (20, 10, 14) {real, imag} */,
  {32'hc18b1dde, 32'hc2772c26} /* (20, 10, 13) {real, imag} */,
  {32'hc07dcb20, 32'h428a53fc} /* (20, 10, 12) {real, imag} */,
  {32'hc2d4a402, 32'hc2ada9ee} /* (20, 10, 11) {real, imag} */,
  {32'h42390a8c, 32'hc2a01aaa} /* (20, 10, 10) {real, imag} */,
  {32'h42baee3c, 32'h40967da8} /* (20, 10, 9) {real, imag} */,
  {32'h42d08b1c, 32'h42257c50} /* (20, 10, 8) {real, imag} */,
  {32'hc1cd4bc0, 32'hc2c0aaf4} /* (20, 10, 7) {real, imag} */,
  {32'h41ff8bcc, 32'h4254fb56} /* (20, 10, 6) {real, imag} */,
  {32'h413c4280, 32'h4215abc0} /* (20, 10, 5) {real, imag} */,
  {32'h42e60bcb, 32'h423d6c0c} /* (20, 10, 4) {real, imag} */,
  {32'hc1ca43ee, 32'h42da1272} /* (20, 10, 3) {real, imag} */,
  {32'h435d4704, 32'h43644b56} /* (20, 10, 2) {real, imag} */,
  {32'hc450a6b0, 32'hc42fe9bc} /* (20, 10, 1) {real, imag} */,
  {32'hc458451b, 32'h00000000} /* (20, 10, 0) {real, imag} */,
  {32'hc50a67a4, 32'h4486fd42} /* (20, 9, 31) {real, imag} */,
  {32'h444f2eae, 32'hc392eb16} /* (20, 9, 30) {real, imag} */,
  {32'hc2388fb0, 32'h41cfa560} /* (20, 9, 29) {real, imag} */,
  {32'hc2811694, 32'h416d2b08} /* (20, 9, 28) {real, imag} */,
  {32'h42dbb7a6, 32'hc2c5720e} /* (20, 9, 27) {real, imag} */,
  {32'hc2b3d220, 32'hc2060945} /* (20, 9, 26) {real, imag} */,
  {32'hc25b022a, 32'h428db748} /* (20, 9, 25) {real, imag} */,
  {32'hc12cc968, 32'hc29f2ae8} /* (20, 9, 24) {real, imag} */,
  {32'h4264cf3b, 32'h428471c0} /* (20, 9, 23) {real, imag} */,
  {32'h41b34898, 32'hc024c848} /* (20, 9, 22) {real, imag} */,
  {32'h41684ada, 32'hc23f15e2} /* (20, 9, 21) {real, imag} */,
  {32'hc2ae036f, 32'hc1099078} /* (20, 9, 20) {real, imag} */,
  {32'h414b21eb, 32'hc1f16c44} /* (20, 9, 19) {real, imag} */,
  {32'h4214c82c, 32'hc1c334fe} /* (20, 9, 18) {real, imag} */,
  {32'hc28548b6, 32'hc1cd570c} /* (20, 9, 17) {real, imag} */,
  {32'h41e3b080, 32'h00000000} /* (20, 9, 16) {real, imag} */,
  {32'hc28548b6, 32'h41cd570c} /* (20, 9, 15) {real, imag} */,
  {32'h4214c82c, 32'h41c334fe} /* (20, 9, 14) {real, imag} */,
  {32'h414b21eb, 32'h41f16c44} /* (20, 9, 13) {real, imag} */,
  {32'hc2ae036f, 32'h41099078} /* (20, 9, 12) {real, imag} */,
  {32'h41684ada, 32'h423f15e2} /* (20, 9, 11) {real, imag} */,
  {32'h41b34898, 32'h4024c848} /* (20, 9, 10) {real, imag} */,
  {32'h4264cf3b, 32'hc28471c0} /* (20, 9, 9) {real, imag} */,
  {32'hc12cc968, 32'h429f2ae8} /* (20, 9, 8) {real, imag} */,
  {32'hc25b022a, 32'hc28db748} /* (20, 9, 7) {real, imag} */,
  {32'hc2b3d220, 32'h42060945} /* (20, 9, 6) {real, imag} */,
  {32'h42dbb7a6, 32'h42c5720e} /* (20, 9, 5) {real, imag} */,
  {32'hc2811694, 32'hc16d2b08} /* (20, 9, 4) {real, imag} */,
  {32'hc2388fb0, 32'hc1cfa560} /* (20, 9, 3) {real, imag} */,
  {32'h444f2eae, 32'h4392eb16} /* (20, 9, 2) {real, imag} */,
  {32'hc50a67a4, 32'hc486fd42} /* (20, 9, 1) {real, imag} */,
  {32'hc50729cd, 32'h00000000} /* (20, 9, 0) {real, imag} */,
  {32'hc5457701, 32'h44c9462d} /* (20, 8, 31) {real, imag} */,
  {32'h4485fa8a, 32'hc3f96f7d} /* (20, 8, 30) {real, imag} */,
  {32'hc2e0086d, 32'h42032dfb} /* (20, 8, 29) {real, imag} */,
  {32'hc20ddfa4, 32'h419a4069} /* (20, 8, 28) {real, imag} */,
  {32'h42f34682, 32'hc1aa3f1c} /* (20, 8, 27) {real, imag} */,
  {32'hc2e53e34, 32'hc2f07234} /* (20, 8, 26) {real, imag} */,
  {32'h41a48fc5, 32'h435986b6} /* (20, 8, 25) {real, imag} */,
  {32'h41aa812b, 32'hc33924e4} /* (20, 8, 24) {real, imag} */,
  {32'hc2961d33, 32'hc24e9ae1} /* (20, 8, 23) {real, imag} */,
  {32'hc29744d6, 32'h4199f18a} /* (20, 8, 22) {real, imag} */,
  {32'hc1897519, 32'hc1c10eb2} /* (20, 8, 21) {real, imag} */,
  {32'h41c3820e, 32'hc1ad55e0} /* (20, 8, 20) {real, imag} */,
  {32'h42d295d3, 32'hc14a71b8} /* (20, 8, 19) {real, imag} */,
  {32'h41d1a4de, 32'hc1c39e23} /* (20, 8, 18) {real, imag} */,
  {32'h41ccb20d, 32'h4269f571} /* (20, 8, 17) {real, imag} */,
  {32'hc1c481e3, 32'h00000000} /* (20, 8, 16) {real, imag} */,
  {32'h41ccb20d, 32'hc269f571} /* (20, 8, 15) {real, imag} */,
  {32'h41d1a4de, 32'h41c39e23} /* (20, 8, 14) {real, imag} */,
  {32'h42d295d3, 32'h414a71b8} /* (20, 8, 13) {real, imag} */,
  {32'h41c3820e, 32'h41ad55e0} /* (20, 8, 12) {real, imag} */,
  {32'hc1897519, 32'h41c10eb2} /* (20, 8, 11) {real, imag} */,
  {32'hc29744d6, 32'hc199f18a} /* (20, 8, 10) {real, imag} */,
  {32'hc2961d33, 32'h424e9ae1} /* (20, 8, 9) {real, imag} */,
  {32'h41aa812b, 32'h433924e4} /* (20, 8, 8) {real, imag} */,
  {32'h41a48fc5, 32'hc35986b6} /* (20, 8, 7) {real, imag} */,
  {32'hc2e53e34, 32'h42f07234} /* (20, 8, 6) {real, imag} */,
  {32'h42f34682, 32'h41aa3f1c} /* (20, 8, 5) {real, imag} */,
  {32'hc20ddfa4, 32'hc19a4069} /* (20, 8, 4) {real, imag} */,
  {32'hc2e0086d, 32'hc2032dfb} /* (20, 8, 3) {real, imag} */,
  {32'h4485fa8a, 32'h43f96f7d} /* (20, 8, 2) {real, imag} */,
  {32'hc5457701, 32'hc4c9462d} /* (20, 8, 1) {real, imag} */,
  {32'hc546e5c6, 32'h00000000} /* (20, 8, 0) {real, imag} */,
  {32'hc56b697f, 32'h44f8227e} /* (20, 7, 31) {real, imag} */,
  {32'h4480347d, 32'hc40eb10b} /* (20, 7, 30) {real, imag} */,
  {32'hc1a05e9c, 32'hc30cdef6} /* (20, 7, 29) {real, imag} */,
  {32'hc2268188, 32'h4256f456} /* (20, 7, 28) {real, imag} */,
  {32'h43846a0c, 32'hc1fe4da0} /* (20, 7, 27) {real, imag} */,
  {32'h41c0f902, 32'hc28534a6} /* (20, 7, 26) {real, imag} */,
  {32'h41d7e577, 32'h427abad1} /* (20, 7, 25) {real, imag} */,
  {32'h42be31a2, 32'hc32d64b0} /* (20, 7, 24) {real, imag} */,
  {32'hc2821945, 32'h422206cf} /* (20, 7, 23) {real, imag} */,
  {32'h41c9fcdb, 32'hc21de380} /* (20, 7, 22) {real, imag} */,
  {32'h4177a620, 32'hc1db8a27} /* (20, 7, 21) {real, imag} */,
  {32'hc2175042, 32'h42d26283} /* (20, 7, 20) {real, imag} */,
  {32'h41a22f7a, 32'hc2603e52} /* (20, 7, 19) {real, imag} */,
  {32'hc17bb2fe, 32'h42573d9f} /* (20, 7, 18) {real, imag} */,
  {32'h41560274, 32'hc2be3158} /* (20, 7, 17) {real, imag} */,
  {32'h3fc7b2b0, 32'h00000000} /* (20, 7, 16) {real, imag} */,
  {32'h41560274, 32'h42be3158} /* (20, 7, 15) {real, imag} */,
  {32'hc17bb2fe, 32'hc2573d9f} /* (20, 7, 14) {real, imag} */,
  {32'h41a22f7a, 32'h42603e52} /* (20, 7, 13) {real, imag} */,
  {32'hc2175042, 32'hc2d26283} /* (20, 7, 12) {real, imag} */,
  {32'h4177a620, 32'h41db8a27} /* (20, 7, 11) {real, imag} */,
  {32'h41c9fcdb, 32'h421de380} /* (20, 7, 10) {real, imag} */,
  {32'hc2821945, 32'hc22206cf} /* (20, 7, 9) {real, imag} */,
  {32'h42be31a2, 32'h432d64b0} /* (20, 7, 8) {real, imag} */,
  {32'h41d7e577, 32'hc27abad1} /* (20, 7, 7) {real, imag} */,
  {32'h41c0f902, 32'h428534a6} /* (20, 7, 6) {real, imag} */,
  {32'h43846a0c, 32'h41fe4da0} /* (20, 7, 5) {real, imag} */,
  {32'hc2268188, 32'hc256f456} /* (20, 7, 4) {real, imag} */,
  {32'hc1a05e9c, 32'h430cdef6} /* (20, 7, 3) {real, imag} */,
  {32'h4480347d, 32'h440eb10b} /* (20, 7, 2) {real, imag} */,
  {32'hc56b697f, 32'hc4f8227e} /* (20, 7, 1) {real, imag} */,
  {32'hc5722bee, 32'h00000000} /* (20, 7, 0) {real, imag} */,
  {32'hc5731306, 32'h4519b901} /* (20, 6, 31) {real, imag} */,
  {32'h44491a31, 32'hc42fbd16} /* (20, 6, 30) {real, imag} */,
  {32'h3fb953c0, 32'h424d60a6} /* (20, 6, 29) {real, imag} */,
  {32'hc2276140, 32'hc21b0eae} /* (20, 6, 28) {real, imag} */,
  {32'h4388c814, 32'h41c9e288} /* (20, 6, 27) {real, imag} */,
  {32'h4131ed97, 32'hc15adb68} /* (20, 6, 26) {real, imag} */,
  {32'hc2d196d0, 32'h424d0969} /* (20, 6, 25) {real, imag} */,
  {32'h41010814, 32'hc23f179e} /* (20, 6, 24) {real, imag} */,
  {32'hc2970194, 32'h43016077} /* (20, 6, 23) {real, imag} */,
  {32'h4247c0a1, 32'hc245e77c} /* (20, 6, 22) {real, imag} */,
  {32'h425c3fac, 32'h41cedda3} /* (20, 6, 21) {real, imag} */,
  {32'hc022b080, 32'hc201d7c4} /* (20, 6, 20) {real, imag} */,
  {32'h415ef3fe, 32'hc1fbd42c} /* (20, 6, 19) {real, imag} */,
  {32'h41ae49bc, 32'h42a61262} /* (20, 6, 18) {real, imag} */,
  {32'h4171a82d, 32'h40946e2e} /* (20, 6, 17) {real, imag} */,
  {32'h41aba05b, 32'h00000000} /* (20, 6, 16) {real, imag} */,
  {32'h4171a82d, 32'hc0946e2e} /* (20, 6, 15) {real, imag} */,
  {32'h41ae49bc, 32'hc2a61262} /* (20, 6, 14) {real, imag} */,
  {32'h415ef3fe, 32'h41fbd42c} /* (20, 6, 13) {real, imag} */,
  {32'hc022b080, 32'h4201d7c4} /* (20, 6, 12) {real, imag} */,
  {32'h425c3fac, 32'hc1cedda3} /* (20, 6, 11) {real, imag} */,
  {32'h4247c0a1, 32'h4245e77c} /* (20, 6, 10) {real, imag} */,
  {32'hc2970194, 32'hc3016077} /* (20, 6, 9) {real, imag} */,
  {32'h41010814, 32'h423f179e} /* (20, 6, 8) {real, imag} */,
  {32'hc2d196d0, 32'hc24d0969} /* (20, 6, 7) {real, imag} */,
  {32'h4131ed97, 32'h415adb68} /* (20, 6, 6) {real, imag} */,
  {32'h4388c814, 32'hc1c9e288} /* (20, 6, 5) {real, imag} */,
  {32'hc2276140, 32'h421b0eae} /* (20, 6, 4) {real, imag} */,
  {32'h3fb953c0, 32'hc24d60a6} /* (20, 6, 3) {real, imag} */,
  {32'h44491a31, 32'h442fbd16} /* (20, 6, 2) {real, imag} */,
  {32'hc5731306, 32'hc519b901} /* (20, 6, 1) {real, imag} */,
  {32'hc583cbcb, 32'h00000000} /* (20, 6, 0) {real, imag} */,
  {32'hc56bef1d, 32'h4547c3d0} /* (20, 5, 31) {real, imag} */,
  {32'h439f980c, 32'hc4534b44} /* (20, 5, 30) {real, imag} */,
  {32'h426f42fc, 32'hc2b33d12} /* (20, 5, 29) {real, imag} */,
  {32'h42cad0ed, 32'hc338a062} /* (20, 5, 28) {real, imag} */,
  {32'h4355ca3f, 32'h42492eb3} /* (20, 5, 27) {real, imag} */,
  {32'h42b3b76b, 32'h42f31c44} /* (20, 5, 26) {real, imag} */,
  {32'hc213fe08, 32'h4298adda} /* (20, 5, 25) {real, imag} */,
  {32'hbf9e9fa0, 32'hc243b22a} /* (20, 5, 24) {real, imag} */,
  {32'h42398567, 32'h4123132c} /* (20, 5, 23) {real, imag} */,
  {32'hc28b6b36, 32'hc2ced4ca} /* (20, 5, 22) {real, imag} */,
  {32'hc2d50a8a, 32'hc20aba27} /* (20, 5, 21) {real, imag} */,
  {32'hc1c619a6, 32'hc234c726} /* (20, 5, 20) {real, imag} */,
  {32'hc25fa118, 32'h4103692c} /* (20, 5, 19) {real, imag} */,
  {32'h42c63796, 32'hc2929b09} /* (20, 5, 18) {real, imag} */,
  {32'h428d3a97, 32'h41e9014a} /* (20, 5, 17) {real, imag} */,
  {32'h4288c66e, 32'h00000000} /* (20, 5, 16) {real, imag} */,
  {32'h428d3a97, 32'hc1e9014a} /* (20, 5, 15) {real, imag} */,
  {32'h42c63796, 32'h42929b09} /* (20, 5, 14) {real, imag} */,
  {32'hc25fa118, 32'hc103692c} /* (20, 5, 13) {real, imag} */,
  {32'hc1c619a6, 32'h4234c726} /* (20, 5, 12) {real, imag} */,
  {32'hc2d50a8a, 32'h420aba27} /* (20, 5, 11) {real, imag} */,
  {32'hc28b6b36, 32'h42ced4ca} /* (20, 5, 10) {real, imag} */,
  {32'h42398567, 32'hc123132c} /* (20, 5, 9) {real, imag} */,
  {32'hbf9e9fa0, 32'h4243b22a} /* (20, 5, 8) {real, imag} */,
  {32'hc213fe08, 32'hc298adda} /* (20, 5, 7) {real, imag} */,
  {32'h42b3b76b, 32'hc2f31c44} /* (20, 5, 6) {real, imag} */,
  {32'h4355ca3f, 32'hc2492eb3} /* (20, 5, 5) {real, imag} */,
  {32'h42cad0ed, 32'h4338a062} /* (20, 5, 4) {real, imag} */,
  {32'h426f42fc, 32'h42b33d12} /* (20, 5, 3) {real, imag} */,
  {32'h439f980c, 32'h44534b44} /* (20, 5, 2) {real, imag} */,
  {32'hc56bef1d, 32'hc547c3d0} /* (20, 5, 1) {real, imag} */,
  {32'hc59025f4, 32'h00000000} /* (20, 5, 0) {real, imag} */,
  {32'hc55d4e0c, 32'h45702e38} /* (20, 4, 31) {real, imag} */,
  {32'hc328390c, 32'hc47a9df2} /* (20, 4, 30) {real, imag} */,
  {32'h428dea14, 32'hc371b47e} /* (20, 4, 29) {real, imag} */,
  {32'h433e78fa, 32'hc3672ae0} /* (20, 4, 28) {real, imag} */,
  {32'h4355dc6d, 32'h4349b2fb} /* (20, 4, 27) {real, imag} */,
  {32'h4100f3ac, 32'h42091ec1} /* (20, 4, 26) {real, imag} */,
  {32'hc211c25c, 32'hc27c704c} /* (20, 4, 25) {real, imag} */,
  {32'hc1b27c96, 32'h416385f4} /* (20, 4, 24) {real, imag} */,
  {32'h42429e4c, 32'h40d65c68} /* (20, 4, 23) {real, imag} */,
  {32'h410fc822, 32'h42667c27} /* (20, 4, 22) {real, imag} */,
  {32'hc22eba4a, 32'hc27b80a6} /* (20, 4, 21) {real, imag} */,
  {32'hc098db7a, 32'h4168df97} /* (20, 4, 20) {real, imag} */,
  {32'hc25380c1, 32'h428a3ae8} /* (20, 4, 19) {real, imag} */,
  {32'hc197768e, 32'hc11e2b4f} /* (20, 4, 18) {real, imag} */,
  {32'hc0065c18, 32'hc2c6ec80} /* (20, 4, 17) {real, imag} */,
  {32'hc1e9c3f7, 32'h00000000} /* (20, 4, 16) {real, imag} */,
  {32'hc0065c18, 32'h42c6ec80} /* (20, 4, 15) {real, imag} */,
  {32'hc197768e, 32'h411e2b4f} /* (20, 4, 14) {real, imag} */,
  {32'hc25380c1, 32'hc28a3ae8} /* (20, 4, 13) {real, imag} */,
  {32'hc098db7a, 32'hc168df97} /* (20, 4, 12) {real, imag} */,
  {32'hc22eba4a, 32'h427b80a6} /* (20, 4, 11) {real, imag} */,
  {32'h410fc822, 32'hc2667c27} /* (20, 4, 10) {real, imag} */,
  {32'h42429e4c, 32'hc0d65c68} /* (20, 4, 9) {real, imag} */,
  {32'hc1b27c96, 32'hc16385f4} /* (20, 4, 8) {real, imag} */,
  {32'hc211c25c, 32'h427c704c} /* (20, 4, 7) {real, imag} */,
  {32'h4100f3ac, 32'hc2091ec1} /* (20, 4, 6) {real, imag} */,
  {32'h4355dc6d, 32'hc349b2fb} /* (20, 4, 5) {real, imag} */,
  {32'h433e78fa, 32'h43672ae0} /* (20, 4, 4) {real, imag} */,
  {32'h428dea14, 32'h4371b47e} /* (20, 4, 3) {real, imag} */,
  {32'hc328390c, 32'h447a9df2} /* (20, 4, 2) {real, imag} */,
  {32'hc55d4e0c, 32'hc5702e38} /* (20, 4, 1) {real, imag} */,
  {32'hc5987be6, 32'h00000000} /* (20, 4, 0) {real, imag} */,
  {32'hc550db8a, 32'h457e9913} /* (20, 3, 31) {real, imag} */,
  {32'hc3dad868, 32'hc49a8313} /* (20, 3, 30) {real, imag} */,
  {32'h410c7c64, 32'hc344e81e} /* (20, 3, 29) {real, imag} */,
  {32'h431eebfa, 32'hc38599a8} /* (20, 3, 28) {real, imag} */,
  {32'h433e6040, 32'h43189d2c} /* (20, 3, 27) {real, imag} */,
  {32'h41b81ca4, 32'h4204635c} /* (20, 3, 26) {real, imag} */,
  {32'h42744e7a, 32'hc277f352} /* (20, 3, 25) {real, imag} */,
  {32'hc21c3924, 32'hc2fa2f7e} /* (20, 3, 24) {real, imag} */,
  {32'h42526489, 32'hc1219b44} /* (20, 3, 23) {real, imag} */,
  {32'h429f378b, 32'hc2dd16d0} /* (20, 3, 22) {real, imag} */,
  {32'h424ec8c2, 32'h42ce0f99} /* (20, 3, 21) {real, imag} */,
  {32'hc2a24422, 32'h41f24e59} /* (20, 3, 20) {real, imag} */,
  {32'hc1432283, 32'hc20dc37c} /* (20, 3, 19) {real, imag} */,
  {32'h42ac780b, 32'hc1940c43} /* (20, 3, 18) {real, imag} */,
  {32'h4285b589, 32'hc19f38a2} /* (20, 3, 17) {real, imag} */,
  {32'h4117d4f8, 32'h00000000} /* (20, 3, 16) {real, imag} */,
  {32'h4285b589, 32'h419f38a2} /* (20, 3, 15) {real, imag} */,
  {32'h42ac780b, 32'h41940c43} /* (20, 3, 14) {real, imag} */,
  {32'hc1432283, 32'h420dc37c} /* (20, 3, 13) {real, imag} */,
  {32'hc2a24422, 32'hc1f24e59} /* (20, 3, 12) {real, imag} */,
  {32'h424ec8c2, 32'hc2ce0f99} /* (20, 3, 11) {real, imag} */,
  {32'h429f378b, 32'h42dd16d0} /* (20, 3, 10) {real, imag} */,
  {32'h42526489, 32'h41219b44} /* (20, 3, 9) {real, imag} */,
  {32'hc21c3924, 32'h42fa2f7e} /* (20, 3, 8) {real, imag} */,
  {32'h42744e7a, 32'h4277f352} /* (20, 3, 7) {real, imag} */,
  {32'h41b81ca4, 32'hc204635c} /* (20, 3, 6) {real, imag} */,
  {32'h433e6040, 32'hc3189d2c} /* (20, 3, 5) {real, imag} */,
  {32'h431eebfa, 32'h438599a8} /* (20, 3, 4) {real, imag} */,
  {32'h410c7c64, 32'h4344e81e} /* (20, 3, 3) {real, imag} */,
  {32'hc3dad868, 32'h449a8313} /* (20, 3, 2) {real, imag} */,
  {32'hc550db8a, 32'hc57e9913} /* (20, 3, 1) {real, imag} */,
  {32'hc5a3e2b8, 32'h00000000} /* (20, 3, 0) {real, imag} */,
  {32'hc553ed5d, 32'h4576213e} /* (20, 2, 31) {real, imag} */,
  {32'hc377fe48, 32'hc48785f2} /* (20, 2, 30) {real, imag} */,
  {32'h42472c89, 32'hc2b6aa2e} /* (20, 2, 29) {real, imag} */,
  {32'h42858166, 32'hc38f8087} /* (20, 2, 28) {real, imag} */,
  {32'h438d556f, 32'h41e2ab3c} /* (20, 2, 27) {real, imag} */,
  {32'h4297aa9c, 32'hc15ddaf6} /* (20, 2, 26) {real, imag} */,
  {32'h41bde348, 32'h4240482c} /* (20, 2, 25) {real, imag} */,
  {32'hc22ce320, 32'h4231d62e} /* (20, 2, 24) {real, imag} */,
  {32'h4246dd62, 32'hc16e4518} /* (20, 2, 23) {real, imag} */,
  {32'hc082d158, 32'hc25c58b4} /* (20, 2, 22) {real, imag} */,
  {32'hbf7dd620, 32'hc089b5d4} /* (20, 2, 21) {real, imag} */,
  {32'hc1c00d12, 32'hc2b87de3} /* (20, 2, 20) {real, imag} */,
  {32'h4207ced8, 32'hc1eb256d} /* (20, 2, 19) {real, imag} */,
  {32'hc236f220, 32'h402127a8} /* (20, 2, 18) {real, imag} */,
  {32'h41e964ad, 32'hc205938e} /* (20, 2, 17) {real, imag} */,
  {32'hc18790d5, 32'h00000000} /* (20, 2, 16) {real, imag} */,
  {32'h41e964ad, 32'h4205938e} /* (20, 2, 15) {real, imag} */,
  {32'hc236f220, 32'hc02127a8} /* (20, 2, 14) {real, imag} */,
  {32'h4207ced8, 32'h41eb256d} /* (20, 2, 13) {real, imag} */,
  {32'hc1c00d12, 32'h42b87de3} /* (20, 2, 12) {real, imag} */,
  {32'hbf7dd620, 32'h4089b5d4} /* (20, 2, 11) {real, imag} */,
  {32'hc082d158, 32'h425c58b4} /* (20, 2, 10) {real, imag} */,
  {32'h4246dd62, 32'h416e4518} /* (20, 2, 9) {real, imag} */,
  {32'hc22ce320, 32'hc231d62e} /* (20, 2, 8) {real, imag} */,
  {32'h41bde348, 32'hc240482c} /* (20, 2, 7) {real, imag} */,
  {32'h4297aa9c, 32'h415ddaf6} /* (20, 2, 6) {real, imag} */,
  {32'h438d556f, 32'hc1e2ab3c} /* (20, 2, 5) {real, imag} */,
  {32'h42858166, 32'h438f8087} /* (20, 2, 4) {real, imag} */,
  {32'h42472c89, 32'h42b6aa2e} /* (20, 2, 3) {real, imag} */,
  {32'hc377fe48, 32'h448785f2} /* (20, 2, 2) {real, imag} */,
  {32'hc553ed5d, 32'hc576213e} /* (20, 2, 1) {real, imag} */,
  {32'hc5aa6a7a, 32'h00000000} /* (20, 2, 0) {real, imag} */,
  {32'hc55d390c, 32'h45625f2e} /* (20, 1, 31) {real, imag} */,
  {32'hc2ee8c68, 32'hc46c5aec} /* (20, 1, 30) {real, imag} */,
  {32'h4325749a, 32'hc2d83578} /* (20, 1, 29) {real, imag} */,
  {32'h4328fe0d, 32'hc38e2907} /* (20, 1, 28) {real, imag} */,
  {32'h434acdaf, 32'h42914d3d} /* (20, 1, 27) {real, imag} */,
  {32'h42ef522a, 32'hc294bb97} /* (20, 1, 26) {real, imag} */,
  {32'hc3067315, 32'h42ad8828} /* (20, 1, 25) {real, imag} */,
  {32'hc2d309d4, 32'h425a6b26} /* (20, 1, 24) {real, imag} */,
  {32'hc29b6558, 32'h42034e92} /* (20, 1, 23) {real, imag} */,
  {32'h422150d3, 32'hc3407668} /* (20, 1, 22) {real, imag} */,
  {32'h42342b10, 32'hc1f71236} /* (20, 1, 21) {real, imag} */,
  {32'h41c6e7e9, 32'h424f215c} /* (20, 1, 20) {real, imag} */,
  {32'hc1344a80, 32'hc201f76b} /* (20, 1, 19) {real, imag} */,
  {32'hc123f567, 32'hc203b192} /* (20, 1, 18) {real, imag} */,
  {32'hc164d20c, 32'hc1c3a13c} /* (20, 1, 17) {real, imag} */,
  {32'hc1910a46, 32'h00000000} /* (20, 1, 16) {real, imag} */,
  {32'hc164d20c, 32'h41c3a13c} /* (20, 1, 15) {real, imag} */,
  {32'hc123f567, 32'h4203b192} /* (20, 1, 14) {real, imag} */,
  {32'hc1344a80, 32'h4201f76b} /* (20, 1, 13) {real, imag} */,
  {32'h41c6e7e9, 32'hc24f215c} /* (20, 1, 12) {real, imag} */,
  {32'h42342b10, 32'h41f71236} /* (20, 1, 11) {real, imag} */,
  {32'h422150d3, 32'h43407668} /* (20, 1, 10) {real, imag} */,
  {32'hc29b6558, 32'hc2034e92} /* (20, 1, 9) {real, imag} */,
  {32'hc2d309d4, 32'hc25a6b26} /* (20, 1, 8) {real, imag} */,
  {32'hc3067315, 32'hc2ad8828} /* (20, 1, 7) {real, imag} */,
  {32'h42ef522a, 32'h4294bb97} /* (20, 1, 6) {real, imag} */,
  {32'h434acdaf, 32'hc2914d3d} /* (20, 1, 5) {real, imag} */,
  {32'h4328fe0d, 32'h438e2907} /* (20, 1, 4) {real, imag} */,
  {32'h4325749a, 32'h42d83578} /* (20, 1, 3) {real, imag} */,
  {32'hc2ee8c68, 32'h446c5aec} /* (20, 1, 2) {real, imag} */,
  {32'hc55d390c, 32'hc5625f2e} /* (20, 1, 1) {real, imag} */,
  {32'hc5a4bfdf, 32'h00000000} /* (20, 1, 0) {real, imag} */,
  {32'hc56a6f8a, 32'h453910d2} /* (20, 0, 31) {real, imag} */,
  {32'h43315638, 32'hc4369ede} /* (20, 0, 30) {real, imag} */,
  {32'h430c328b, 32'hc1692694} /* (20, 0, 29) {real, imag} */,
  {32'h42047b80, 32'hc318d99e} /* (20, 0, 28) {real, imag} */,
  {32'h41c53dd0, 32'hc0623b10} /* (20, 0, 27) {real, imag} */,
  {32'hc1fcc9b7, 32'hc28ef007} /* (20, 0, 26) {real, imag} */,
  {32'hc29577b1, 32'h418a0036} /* (20, 0, 25) {real, imag} */,
  {32'hc1aaf2f5, 32'hc28e997e} /* (20, 0, 24) {real, imag} */,
  {32'hc23a59d1, 32'h4283b693} /* (20, 0, 23) {real, imag} */,
  {32'hc22b648c, 32'hc2a171f0} /* (20, 0, 22) {real, imag} */,
  {32'h415d1d58, 32'hc070d738} /* (20, 0, 21) {real, imag} */,
  {32'hc1acd2ce, 32'hc234cff2} /* (20, 0, 20) {real, imag} */,
  {32'hc228b89e, 32'hc1a22f96} /* (20, 0, 19) {real, imag} */,
  {32'hc2685a26, 32'hc2192bb5} /* (20, 0, 18) {real, imag} */,
  {32'hc1ee4ed3, 32'h41650b3c} /* (20, 0, 17) {real, imag} */,
  {32'hc184a64c, 32'h00000000} /* (20, 0, 16) {real, imag} */,
  {32'hc1ee4ed3, 32'hc1650b3c} /* (20, 0, 15) {real, imag} */,
  {32'hc2685a26, 32'h42192bb5} /* (20, 0, 14) {real, imag} */,
  {32'hc228b89e, 32'h41a22f96} /* (20, 0, 13) {real, imag} */,
  {32'hc1acd2ce, 32'h4234cff2} /* (20, 0, 12) {real, imag} */,
  {32'h415d1d58, 32'h4070d738} /* (20, 0, 11) {real, imag} */,
  {32'hc22b648c, 32'h42a171f0} /* (20, 0, 10) {real, imag} */,
  {32'hc23a59d1, 32'hc283b693} /* (20, 0, 9) {real, imag} */,
  {32'hc1aaf2f5, 32'h428e997e} /* (20, 0, 8) {real, imag} */,
  {32'hc29577b1, 32'hc18a0036} /* (20, 0, 7) {real, imag} */,
  {32'hc1fcc9b7, 32'h428ef007} /* (20, 0, 6) {real, imag} */,
  {32'h41c53dd0, 32'h40623b10} /* (20, 0, 5) {real, imag} */,
  {32'h42047b80, 32'h4318d99e} /* (20, 0, 4) {real, imag} */,
  {32'h430c328b, 32'h41692694} /* (20, 0, 3) {real, imag} */,
  {32'h43315638, 32'h44369ede} /* (20, 0, 2) {real, imag} */,
  {32'hc56a6f8a, 32'hc53910d2} /* (20, 0, 1) {real, imag} */,
  {32'hc59efb64, 32'h00000000} /* (20, 0, 0) {real, imag} */,
  {32'hc576fb87, 32'h44fd39e8} /* (19, 31, 31) {real, imag} */,
  {32'h44235dba, 32'hc3fed87d} /* (19, 31, 30) {real, imag} */,
  {32'h423032f2, 32'h41c0572a} /* (19, 31, 29) {real, imag} */,
  {32'hc201ffe9, 32'h3fca6b80} /* (19, 31, 28) {real, imag} */,
  {32'h429795c1, 32'hc29b7899} /* (19, 31, 27) {real, imag} */,
  {32'hc248693c, 32'h41b15064} /* (19, 31, 26) {real, imag} */,
  {32'hc2280d40, 32'h41758820} /* (19, 31, 25) {real, imag} */,
  {32'h4296b18f, 32'hc232f5a6} /* (19, 31, 24) {real, imag} */,
  {32'h42ddb5b3, 32'h41eaf9fc} /* (19, 31, 23) {real, imag} */,
  {32'h419efee7, 32'hc29edebf} /* (19, 31, 22) {real, imag} */,
  {32'h426851c8, 32'h418f2d9c} /* (19, 31, 21) {real, imag} */,
  {32'hc18dcab0, 32'hc11ce8da} /* (19, 31, 20) {real, imag} */,
  {32'hc1e392f8, 32'hc19cdabd} /* (19, 31, 19) {real, imag} */,
  {32'h40a14828, 32'hc1896951} /* (19, 31, 18) {real, imag} */,
  {32'hc1816777, 32'h40d11074} /* (19, 31, 17) {real, imag} */,
  {32'hc23b2661, 32'h00000000} /* (19, 31, 16) {real, imag} */,
  {32'hc1816777, 32'hc0d11074} /* (19, 31, 15) {real, imag} */,
  {32'h40a14828, 32'h41896951} /* (19, 31, 14) {real, imag} */,
  {32'hc1e392f8, 32'h419cdabd} /* (19, 31, 13) {real, imag} */,
  {32'hc18dcab0, 32'h411ce8da} /* (19, 31, 12) {real, imag} */,
  {32'h426851c8, 32'hc18f2d9c} /* (19, 31, 11) {real, imag} */,
  {32'h419efee7, 32'h429edebf} /* (19, 31, 10) {real, imag} */,
  {32'h42ddb5b3, 32'hc1eaf9fc} /* (19, 31, 9) {real, imag} */,
  {32'h4296b18f, 32'h4232f5a6} /* (19, 31, 8) {real, imag} */,
  {32'hc2280d40, 32'hc1758820} /* (19, 31, 7) {real, imag} */,
  {32'hc248693c, 32'hc1b15064} /* (19, 31, 6) {real, imag} */,
  {32'h429795c1, 32'h429b7899} /* (19, 31, 5) {real, imag} */,
  {32'hc201ffe9, 32'hbfca6b80} /* (19, 31, 4) {real, imag} */,
  {32'h423032f2, 32'hc1c0572a} /* (19, 31, 3) {real, imag} */,
  {32'h44235dba, 32'h43fed87d} /* (19, 31, 2) {real, imag} */,
  {32'hc576fb87, 32'hc4fd39e8} /* (19, 31, 1) {real, imag} */,
  {32'hc594785b, 32'h00000000} /* (19, 31, 0) {real, imag} */,
  {32'hc58d91ce, 32'h44d6ba0c} /* (19, 30, 31) {real, imag} */,
  {32'h449936ee, 32'hc3f272f4} /* (19, 30, 30) {real, imag} */,
  {32'h4251c236, 32'hc10d1b50} /* (19, 30, 29) {real, imag} */,
  {32'hc246236b, 32'h42129818} /* (19, 30, 28) {real, imag} */,
  {32'h423fc38e, 32'hc2cb0d84} /* (19, 30, 27) {real, imag} */,
  {32'h423d58ce, 32'h404ad480} /* (19, 30, 26) {real, imag} */,
  {32'h420fffa4, 32'h42ff5508} /* (19, 30, 25) {real, imag} */,
  {32'h427381e2, 32'h413a42d8} /* (19, 30, 24) {real, imag} */,
  {32'h42a6e160, 32'hc2ee0cc0} /* (19, 30, 23) {real, imag} */,
  {32'h40d38d48, 32'hc25342a8} /* (19, 30, 22) {real, imag} */,
  {32'hc2830a84, 32'hc283f030} /* (19, 30, 21) {real, imag} */,
  {32'h41b7d902, 32'h421de7ba} /* (19, 30, 20) {real, imag} */,
  {32'h422b92cb, 32'h423bbcc8} /* (19, 30, 19) {real, imag} */,
  {32'hc0b2534f, 32'hc26e35e2} /* (19, 30, 18) {real, imag} */,
  {32'hc26271ee, 32'hc226eed3} /* (19, 30, 17) {real, imag} */,
  {32'h42645f63, 32'h00000000} /* (19, 30, 16) {real, imag} */,
  {32'hc26271ee, 32'h4226eed3} /* (19, 30, 15) {real, imag} */,
  {32'hc0b2534f, 32'h426e35e2} /* (19, 30, 14) {real, imag} */,
  {32'h422b92cb, 32'hc23bbcc8} /* (19, 30, 13) {real, imag} */,
  {32'h41b7d902, 32'hc21de7ba} /* (19, 30, 12) {real, imag} */,
  {32'hc2830a84, 32'h4283f030} /* (19, 30, 11) {real, imag} */,
  {32'h40d38d48, 32'h425342a8} /* (19, 30, 10) {real, imag} */,
  {32'h42a6e160, 32'h42ee0cc0} /* (19, 30, 9) {real, imag} */,
  {32'h427381e2, 32'hc13a42d8} /* (19, 30, 8) {real, imag} */,
  {32'h420fffa4, 32'hc2ff5508} /* (19, 30, 7) {real, imag} */,
  {32'h423d58ce, 32'hc04ad480} /* (19, 30, 6) {real, imag} */,
  {32'h423fc38e, 32'h42cb0d84} /* (19, 30, 5) {real, imag} */,
  {32'hc246236b, 32'hc2129818} /* (19, 30, 4) {real, imag} */,
  {32'h4251c236, 32'h410d1b50} /* (19, 30, 3) {real, imag} */,
  {32'h449936ee, 32'h43f272f4} /* (19, 30, 2) {real, imag} */,
  {32'hc58d91ce, 32'hc4d6ba0c} /* (19, 30, 1) {real, imag} */,
  {32'hc59707b5, 32'h00000000} /* (19, 30, 0) {real, imag} */,
  {32'hc5969d16, 32'h44a75245} /* (19, 29, 31) {real, imag} */,
  {32'h44b89a72, 32'hc3ebdd98} /* (19, 29, 30) {real, imag} */,
  {32'h412fd496, 32'hc296a6ad} /* (19, 29, 29) {real, imag} */,
  {32'hc3a47189, 32'h42c918a1} /* (19, 29, 28) {real, imag} */,
  {32'h432182b2, 32'hc19b1388} /* (19, 29, 27) {real, imag} */,
  {32'h41ca54ee, 32'hc2aba309} /* (19, 29, 26) {real, imag} */,
  {32'hc28c0232, 32'hc10b829c} /* (19, 29, 25) {real, imag} */,
  {32'h3fae3990, 32'h42d1a966} /* (19, 29, 24) {real, imag} */,
  {32'h41bd2fc0, 32'hc2e6f89a} /* (19, 29, 23) {real, imag} */,
  {32'hc16b0c09, 32'h426d1528} /* (19, 29, 22) {real, imag} */,
  {32'h42310686, 32'hc101744a} /* (19, 29, 21) {real, imag} */,
  {32'hc217af6d, 32'h413fdb36} /* (19, 29, 20) {real, imag} */,
  {32'h4234bfdf, 32'h40feda38} /* (19, 29, 19) {real, imag} */,
  {32'h41371b3c, 32'hc2a9bcd5} /* (19, 29, 18) {real, imag} */,
  {32'h3fbe5ff8, 32'h405b9ffe} /* (19, 29, 17) {real, imag} */,
  {32'h42bb2db0, 32'h00000000} /* (19, 29, 16) {real, imag} */,
  {32'h3fbe5ff8, 32'hc05b9ffe} /* (19, 29, 15) {real, imag} */,
  {32'h41371b3c, 32'h42a9bcd5} /* (19, 29, 14) {real, imag} */,
  {32'h4234bfdf, 32'hc0feda38} /* (19, 29, 13) {real, imag} */,
  {32'hc217af6d, 32'hc13fdb36} /* (19, 29, 12) {real, imag} */,
  {32'h42310686, 32'h4101744a} /* (19, 29, 11) {real, imag} */,
  {32'hc16b0c09, 32'hc26d1528} /* (19, 29, 10) {real, imag} */,
  {32'h41bd2fc0, 32'h42e6f89a} /* (19, 29, 9) {real, imag} */,
  {32'h3fae3990, 32'hc2d1a966} /* (19, 29, 8) {real, imag} */,
  {32'hc28c0232, 32'h410b829c} /* (19, 29, 7) {real, imag} */,
  {32'h41ca54ee, 32'h42aba309} /* (19, 29, 6) {real, imag} */,
  {32'h432182b2, 32'h419b1388} /* (19, 29, 5) {real, imag} */,
  {32'hc3a47189, 32'hc2c918a1} /* (19, 29, 4) {real, imag} */,
  {32'h412fd496, 32'h4296a6ad} /* (19, 29, 3) {real, imag} */,
  {32'h44b89a72, 32'h43ebdd98} /* (19, 29, 2) {real, imag} */,
  {32'hc5969d16, 32'hc4a75245} /* (19, 29, 1) {real, imag} */,
  {32'hc595f1d5, 32'h00000000} /* (19, 29, 0) {real, imag} */,
  {32'hc59cd23a, 32'h449d2dcf} /* (19, 28, 31) {real, imag} */,
  {32'h44cf83f8, 32'hc3a4066c} /* (19, 28, 30) {real, imag} */,
  {32'h41ebe6e6, 32'hc333cdba} /* (19, 28, 29) {real, imag} */,
  {32'hc39608c0, 32'h427e7fd6} /* (19, 28, 28) {real, imag} */,
  {32'h4347af47, 32'hbe994200} /* (19, 28, 27) {real, imag} */,
  {32'h42988034, 32'hc2f8e296} /* (19, 28, 26) {real, imag} */,
  {32'hc2a877dc, 32'hc2b819ea} /* (19, 28, 25) {real, imag} */,
  {32'hbfa09d50, 32'hc2041b71} /* (19, 28, 24) {real, imag} */,
  {32'hc2883e3e, 32'h3fbfb7d8} /* (19, 28, 23) {real, imag} */,
  {32'h42322218, 32'h42cc7918} /* (19, 28, 22) {real, imag} */,
  {32'h41006e20, 32'hc252978a} /* (19, 28, 21) {real, imag} */,
  {32'hc1a0a315, 32'hc1f398f6} /* (19, 28, 20) {real, imag} */,
  {32'h426fcc85, 32'h42934809} /* (19, 28, 19) {real, imag} */,
  {32'h42edca07, 32'hc2fb67d1} /* (19, 28, 18) {real, imag} */,
  {32'hc29f1e07, 32'hc188494b} /* (19, 28, 17) {real, imag} */,
  {32'hc1db10e0, 32'h00000000} /* (19, 28, 16) {real, imag} */,
  {32'hc29f1e07, 32'h4188494b} /* (19, 28, 15) {real, imag} */,
  {32'h42edca07, 32'h42fb67d1} /* (19, 28, 14) {real, imag} */,
  {32'h426fcc85, 32'hc2934809} /* (19, 28, 13) {real, imag} */,
  {32'hc1a0a315, 32'h41f398f6} /* (19, 28, 12) {real, imag} */,
  {32'h41006e20, 32'h4252978a} /* (19, 28, 11) {real, imag} */,
  {32'h42322218, 32'hc2cc7918} /* (19, 28, 10) {real, imag} */,
  {32'hc2883e3e, 32'hbfbfb7d8} /* (19, 28, 9) {real, imag} */,
  {32'hbfa09d50, 32'h42041b71} /* (19, 28, 8) {real, imag} */,
  {32'hc2a877dc, 32'h42b819ea} /* (19, 28, 7) {real, imag} */,
  {32'h42988034, 32'h42f8e296} /* (19, 28, 6) {real, imag} */,
  {32'h4347af47, 32'h3e994200} /* (19, 28, 5) {real, imag} */,
  {32'hc39608c0, 32'hc27e7fd6} /* (19, 28, 4) {real, imag} */,
  {32'h41ebe6e6, 32'h4333cdba} /* (19, 28, 3) {real, imag} */,
  {32'h44cf83f8, 32'h43a4066c} /* (19, 28, 2) {real, imag} */,
  {32'hc59cd23a, 32'hc49d2dcf} /* (19, 28, 1) {real, imag} */,
  {32'hc599e26a, 32'h00000000} /* (19, 28, 0) {real, imag} */,
  {32'hc5991ac2, 32'h446c0b70} /* (19, 27, 31) {real, imag} */,
  {32'h44debbac, 32'hc3cef1f0} /* (19, 27, 30) {real, imag} */,
  {32'hc20b9763, 32'hc169ace8} /* (19, 27, 29) {real, imag} */,
  {32'hc38e6ecb, 32'h4135ea90} /* (19, 27, 28) {real, imag} */,
  {32'h42dd4d7a, 32'h4317a038} /* (19, 27, 27) {real, imag} */,
  {32'h42c451c0, 32'h428495f7} /* (19, 27, 26) {real, imag} */,
  {32'hc15b6c50, 32'hc1c1caed} /* (19, 27, 25) {real, imag} */,
  {32'h41bc78ea, 32'hc3128311} /* (19, 27, 24) {real, imag} */,
  {32'h40fe6eb4, 32'hc19dcc48} /* (19, 27, 23) {real, imag} */,
  {32'h41796f34, 32'h425fb0ee} /* (19, 27, 22) {real, imag} */,
  {32'hbf4ddfc0, 32'hc2891f1a} /* (19, 27, 21) {real, imag} */,
  {32'h415de8dd, 32'h3ffc3db0} /* (19, 27, 20) {real, imag} */,
  {32'h42677190, 32'hc21a2f30} /* (19, 27, 19) {real, imag} */,
  {32'hc246abce, 32'h42704386} /* (19, 27, 18) {real, imag} */,
  {32'h4158d24b, 32'h41c72c30} /* (19, 27, 17) {real, imag} */,
  {32'h42ac5172, 32'h00000000} /* (19, 27, 16) {real, imag} */,
  {32'h4158d24b, 32'hc1c72c30} /* (19, 27, 15) {real, imag} */,
  {32'hc246abce, 32'hc2704386} /* (19, 27, 14) {real, imag} */,
  {32'h42677190, 32'h421a2f30} /* (19, 27, 13) {real, imag} */,
  {32'h415de8dd, 32'hbffc3db0} /* (19, 27, 12) {real, imag} */,
  {32'hbf4ddfc0, 32'h42891f1a} /* (19, 27, 11) {real, imag} */,
  {32'h41796f34, 32'hc25fb0ee} /* (19, 27, 10) {real, imag} */,
  {32'h40fe6eb4, 32'h419dcc48} /* (19, 27, 9) {real, imag} */,
  {32'h41bc78ea, 32'h43128311} /* (19, 27, 8) {real, imag} */,
  {32'hc15b6c50, 32'h41c1caed} /* (19, 27, 7) {real, imag} */,
  {32'h42c451c0, 32'hc28495f7} /* (19, 27, 6) {real, imag} */,
  {32'h42dd4d7a, 32'hc317a038} /* (19, 27, 5) {real, imag} */,
  {32'hc38e6ecb, 32'hc135ea90} /* (19, 27, 4) {real, imag} */,
  {32'hc20b9763, 32'h4169ace8} /* (19, 27, 3) {real, imag} */,
  {32'h44debbac, 32'h43cef1f0} /* (19, 27, 2) {real, imag} */,
  {32'hc5991ac2, 32'hc46c0b70} /* (19, 27, 1) {real, imag} */,
  {32'hc59b4138, 32'h00000000} /* (19, 27, 0) {real, imag} */,
  {32'hc5940748, 32'h4442045b} /* (19, 26, 31) {real, imag} */,
  {32'h44d7f53e, 32'hc3f896e5} /* (19, 26, 30) {real, imag} */,
  {32'hc1c4dea4, 32'h4306451c} /* (19, 26, 29) {real, imag} */,
  {32'hc3a1d98a, 32'hc208822b} /* (19, 26, 28) {real, imag} */,
  {32'h4324f27c, 32'hc2b880be} /* (19, 26, 27) {real, imag} */,
  {32'hc1b2ec9e, 32'hc25e16fe} /* (19, 26, 26) {real, imag} */,
  {32'hc22167b4, 32'hc1e274ca} /* (19, 26, 25) {real, imag} */,
  {32'hc2e8023b, 32'hc236536e} /* (19, 26, 24) {real, imag} */,
  {32'h408d5642, 32'hc28ae54d} /* (19, 26, 23) {real, imag} */,
  {32'h41e36c5d, 32'h41efbfc4} /* (19, 26, 22) {real, imag} */,
  {32'h428494c5, 32'h42966074} /* (19, 26, 21) {real, imag} */,
  {32'hc1b87756, 32'hc1e215e0} /* (19, 26, 20) {real, imag} */,
  {32'h42656234, 32'hc289c95e} /* (19, 26, 19) {real, imag} */,
  {32'hc28b7a0d, 32'h3fab6010} /* (19, 26, 18) {real, imag} */,
  {32'h421b94c2, 32'hc0ef8cda} /* (19, 26, 17) {real, imag} */,
  {32'hc1d60978, 32'h00000000} /* (19, 26, 16) {real, imag} */,
  {32'h421b94c2, 32'h40ef8cda} /* (19, 26, 15) {real, imag} */,
  {32'hc28b7a0d, 32'hbfab6010} /* (19, 26, 14) {real, imag} */,
  {32'h42656234, 32'h4289c95e} /* (19, 26, 13) {real, imag} */,
  {32'hc1b87756, 32'h41e215e0} /* (19, 26, 12) {real, imag} */,
  {32'h428494c5, 32'hc2966074} /* (19, 26, 11) {real, imag} */,
  {32'h41e36c5d, 32'hc1efbfc4} /* (19, 26, 10) {real, imag} */,
  {32'h408d5642, 32'h428ae54d} /* (19, 26, 9) {real, imag} */,
  {32'hc2e8023b, 32'h4236536e} /* (19, 26, 8) {real, imag} */,
  {32'hc22167b4, 32'h41e274ca} /* (19, 26, 7) {real, imag} */,
  {32'hc1b2ec9e, 32'h425e16fe} /* (19, 26, 6) {real, imag} */,
  {32'h4324f27c, 32'h42b880be} /* (19, 26, 5) {real, imag} */,
  {32'hc3a1d98a, 32'h4208822b} /* (19, 26, 4) {real, imag} */,
  {32'hc1c4dea4, 32'hc306451c} /* (19, 26, 3) {real, imag} */,
  {32'h44d7f53e, 32'h43f896e5} /* (19, 26, 2) {real, imag} */,
  {32'hc5940748, 32'hc442045b} /* (19, 26, 1) {real, imag} */,
  {32'hc5969ca8, 32'h00000000} /* (19, 26, 0) {real, imag} */,
  {32'hc58bb26a, 32'h442ad46b} /* (19, 25, 31) {real, imag} */,
  {32'h44cf5bda, 32'hc3c1b0a3} /* (19, 25, 30) {real, imag} */,
  {32'hc2a61df6, 32'h41a8de0e} /* (19, 25, 29) {real, imag} */,
  {32'hc3cbb264, 32'hc19e8758} /* (19, 25, 28) {real, imag} */,
  {32'h4383f70c, 32'hc3881acf} /* (19, 25, 27) {real, imag} */,
  {32'hc2f36280, 32'hc27b56f0} /* (19, 25, 26) {real, imag} */,
  {32'h42c5cc90, 32'h42b99f31} /* (19, 25, 25) {real, imag} */,
  {32'h42af53c4, 32'hc211d155} /* (19, 25, 24) {real, imag} */,
  {32'hc1639993, 32'hc331308f} /* (19, 25, 23) {real, imag} */,
  {32'h42b01916, 32'hc0e77b20} /* (19, 25, 22) {real, imag} */,
  {32'h41641110, 32'hc23d9292} /* (19, 25, 21) {real, imag} */,
  {32'h4221107e, 32'hc2550bf8} /* (19, 25, 20) {real, imag} */,
  {32'h429501a9, 32'h425a5452} /* (19, 25, 19) {real, imag} */,
  {32'hc1ffb3e5, 32'hc20f773a} /* (19, 25, 18) {real, imag} */,
  {32'h429102b6, 32'h4206be8c} /* (19, 25, 17) {real, imag} */,
  {32'hc2b26dd6, 32'h00000000} /* (19, 25, 16) {real, imag} */,
  {32'h429102b6, 32'hc206be8c} /* (19, 25, 15) {real, imag} */,
  {32'hc1ffb3e5, 32'h420f773a} /* (19, 25, 14) {real, imag} */,
  {32'h429501a9, 32'hc25a5452} /* (19, 25, 13) {real, imag} */,
  {32'h4221107e, 32'h42550bf8} /* (19, 25, 12) {real, imag} */,
  {32'h41641110, 32'h423d9292} /* (19, 25, 11) {real, imag} */,
  {32'h42b01916, 32'h40e77b20} /* (19, 25, 10) {real, imag} */,
  {32'hc1639993, 32'h4331308f} /* (19, 25, 9) {real, imag} */,
  {32'h42af53c4, 32'h4211d155} /* (19, 25, 8) {real, imag} */,
  {32'h42c5cc90, 32'hc2b99f31} /* (19, 25, 7) {real, imag} */,
  {32'hc2f36280, 32'h427b56f0} /* (19, 25, 6) {real, imag} */,
  {32'h4383f70c, 32'h43881acf} /* (19, 25, 5) {real, imag} */,
  {32'hc3cbb264, 32'h419e8758} /* (19, 25, 4) {real, imag} */,
  {32'hc2a61df6, 32'hc1a8de0e} /* (19, 25, 3) {real, imag} */,
  {32'h44cf5bda, 32'h43c1b0a3} /* (19, 25, 2) {real, imag} */,
  {32'hc58bb26a, 32'hc42ad46b} /* (19, 25, 1) {real, imag} */,
  {32'hc5911c77, 32'h00000000} /* (19, 25, 0) {real, imag} */,
  {32'hc5744cd9, 32'h43bd5e8c} /* (19, 24, 31) {real, imag} */,
  {32'h44d301f9, 32'hc3a1c462} /* (19, 24, 30) {real, imag} */,
  {32'hc312aa6f, 32'hc2496de2} /* (19, 24, 29) {real, imag} */,
  {32'hc3c71592, 32'h40a99510} /* (19, 24, 28) {real, imag} */,
  {32'h43883a66, 32'hc321557e} /* (19, 24, 27) {real, imag} */,
  {32'h423d995b, 32'hc2ea3105} /* (19, 24, 26) {real, imag} */,
  {32'hc293a75a, 32'h42fa6143} /* (19, 24, 25) {real, imag} */,
  {32'hc1032c0c, 32'hc1d05db8} /* (19, 24, 24) {real, imag} */,
  {32'h42fec978, 32'hc1df2cd7} /* (19, 24, 23) {real, imag} */,
  {32'hc1dc4018, 32'hc222f45c} /* (19, 24, 22) {real, imag} */,
  {32'h42855dda, 32'hc0ee1b90} /* (19, 24, 21) {real, imag} */,
  {32'hc192b9a6, 32'h42511000} /* (19, 24, 20) {real, imag} */,
  {32'hc1ca5400, 32'hc297263e} /* (19, 24, 19) {real, imag} */,
  {32'hc227491e, 32'h40936698} /* (19, 24, 18) {real, imag} */,
  {32'hc1fadc4a, 32'h42bf8c9d} /* (19, 24, 17) {real, imag} */,
  {32'h42f62dc0, 32'h00000000} /* (19, 24, 16) {real, imag} */,
  {32'hc1fadc4a, 32'hc2bf8c9d} /* (19, 24, 15) {real, imag} */,
  {32'hc227491e, 32'hc0936698} /* (19, 24, 14) {real, imag} */,
  {32'hc1ca5400, 32'h4297263e} /* (19, 24, 13) {real, imag} */,
  {32'hc192b9a6, 32'hc2511000} /* (19, 24, 12) {real, imag} */,
  {32'h42855dda, 32'h40ee1b90} /* (19, 24, 11) {real, imag} */,
  {32'hc1dc4018, 32'h4222f45c} /* (19, 24, 10) {real, imag} */,
  {32'h42fec978, 32'h41df2cd7} /* (19, 24, 9) {real, imag} */,
  {32'hc1032c0c, 32'h41d05db8} /* (19, 24, 8) {real, imag} */,
  {32'hc293a75a, 32'hc2fa6143} /* (19, 24, 7) {real, imag} */,
  {32'h423d995b, 32'h42ea3105} /* (19, 24, 6) {real, imag} */,
  {32'h43883a66, 32'h4321557e} /* (19, 24, 5) {real, imag} */,
  {32'hc3c71592, 32'hc0a99510} /* (19, 24, 4) {real, imag} */,
  {32'hc312aa6f, 32'h42496de2} /* (19, 24, 3) {real, imag} */,
  {32'h44d301f9, 32'h43a1c462} /* (19, 24, 2) {real, imag} */,
  {32'hc5744cd9, 32'hc3bd5e8c} /* (19, 24, 1) {real, imag} */,
  {32'hc57c1780, 32'h00000000} /* (19, 24, 0) {real, imag} */,
  {32'hc54b8c67, 32'h43a63e90} /* (19, 23, 31) {real, imag} */,
  {32'h44be36c4, 32'hc3b8c0dd} /* (19, 23, 30) {real, imag} */,
  {32'hc341a308, 32'hc33f17ed} /* (19, 23, 29) {real, imag} */,
  {32'hc381432d, 32'h435cd5c3} /* (19, 23, 28) {real, imag} */,
  {32'h43a6a070, 32'hc26778f0} /* (19, 23, 27) {real, imag} */,
  {32'hc2c4806d, 32'hc2a53ddf} /* (19, 23, 26) {real, imag} */,
  {32'hc2495094, 32'h40eb3ed4} /* (19, 23, 25) {real, imag} */,
  {32'h42165742, 32'hc2d6738e} /* (19, 23, 24) {real, imag} */,
  {32'h4293fd33, 32'h42eb9da8} /* (19, 23, 23) {real, imag} */,
  {32'hc1192634, 32'hc22b4f6c} /* (19, 23, 22) {real, imag} */,
  {32'h42b85053, 32'h41947ef0} /* (19, 23, 21) {real, imag} */,
  {32'hbed928a0, 32'h41fefb9b} /* (19, 23, 20) {real, imag} */,
  {32'hc1568e18, 32'hc1faf8b2} /* (19, 23, 19) {real, imag} */,
  {32'h42cda78f, 32'hc24dad15} /* (19, 23, 18) {real, imag} */,
  {32'hc2680bea, 32'h416e1a5e} /* (19, 23, 17) {real, imag} */,
  {32'h4284a396, 32'h00000000} /* (19, 23, 16) {real, imag} */,
  {32'hc2680bea, 32'hc16e1a5e} /* (19, 23, 15) {real, imag} */,
  {32'h42cda78f, 32'h424dad15} /* (19, 23, 14) {real, imag} */,
  {32'hc1568e18, 32'h41faf8b2} /* (19, 23, 13) {real, imag} */,
  {32'hbed928a0, 32'hc1fefb9b} /* (19, 23, 12) {real, imag} */,
  {32'h42b85053, 32'hc1947ef0} /* (19, 23, 11) {real, imag} */,
  {32'hc1192634, 32'h422b4f6c} /* (19, 23, 10) {real, imag} */,
  {32'h4293fd33, 32'hc2eb9da8} /* (19, 23, 9) {real, imag} */,
  {32'h42165742, 32'h42d6738e} /* (19, 23, 8) {real, imag} */,
  {32'hc2495094, 32'hc0eb3ed4} /* (19, 23, 7) {real, imag} */,
  {32'hc2c4806d, 32'h42a53ddf} /* (19, 23, 6) {real, imag} */,
  {32'h43a6a070, 32'h426778f0} /* (19, 23, 5) {real, imag} */,
  {32'hc381432d, 32'hc35cd5c3} /* (19, 23, 4) {real, imag} */,
  {32'hc341a308, 32'h433f17ed} /* (19, 23, 3) {real, imag} */,
  {32'h44be36c4, 32'h43b8c0dd} /* (19, 23, 2) {real, imag} */,
  {32'hc54b8c67, 32'hc3a63e90} /* (19, 23, 1) {real, imag} */,
  {32'hc5566e1a, 32'h00000000} /* (19, 23, 0) {real, imag} */,
  {32'hc511d2e7, 32'h435b2428} /* (19, 22, 31) {real, imag} */,
  {32'h44797bab, 32'hc2fe8bfa} /* (19, 22, 30) {real, imag} */,
  {32'hc339e389, 32'h42983d6e} /* (19, 22, 29) {real, imag} */,
  {32'hc32e2d94, 32'hc1fbb686} /* (19, 22, 28) {real, imag} */,
  {32'h43737156, 32'hc35d73d9} /* (19, 22, 27) {real, imag} */,
  {32'hc21a2ee8, 32'hc2e29fd8} /* (19, 22, 26) {real, imag} */,
  {32'hc22123d4, 32'hc18fcdbe} /* (19, 22, 25) {real, imag} */,
  {32'h42b20b24, 32'hc2813344} /* (19, 22, 24) {real, imag} */,
  {32'hc0bc922c, 32'hc2d7c5ef} /* (19, 22, 23) {real, imag} */,
  {32'h41c2df0e, 32'hc1cc504f} /* (19, 22, 22) {real, imag} */,
  {32'hc28ab78f, 32'hc3164ae4} /* (19, 22, 21) {real, imag} */,
  {32'h42c2fb5a, 32'hc1a83b09} /* (19, 22, 20) {real, imag} */,
  {32'hc20ba668, 32'h42836e55} /* (19, 22, 19) {real, imag} */,
  {32'hc1b42cbc, 32'hc1ecf419} /* (19, 22, 18) {real, imag} */,
  {32'hc24cffb4, 32'h418731c0} /* (19, 22, 17) {real, imag} */,
  {32'hc28cd31a, 32'h00000000} /* (19, 22, 16) {real, imag} */,
  {32'hc24cffb4, 32'hc18731c0} /* (19, 22, 15) {real, imag} */,
  {32'hc1b42cbc, 32'h41ecf419} /* (19, 22, 14) {real, imag} */,
  {32'hc20ba668, 32'hc2836e55} /* (19, 22, 13) {real, imag} */,
  {32'h42c2fb5a, 32'h41a83b09} /* (19, 22, 12) {real, imag} */,
  {32'hc28ab78f, 32'h43164ae4} /* (19, 22, 11) {real, imag} */,
  {32'h41c2df0e, 32'h41cc504f} /* (19, 22, 10) {real, imag} */,
  {32'hc0bc922c, 32'h42d7c5ef} /* (19, 22, 9) {real, imag} */,
  {32'h42b20b24, 32'h42813344} /* (19, 22, 8) {real, imag} */,
  {32'hc22123d4, 32'h418fcdbe} /* (19, 22, 7) {real, imag} */,
  {32'hc21a2ee8, 32'h42e29fd8} /* (19, 22, 6) {real, imag} */,
  {32'h43737156, 32'h435d73d9} /* (19, 22, 5) {real, imag} */,
  {32'hc32e2d94, 32'h41fbb686} /* (19, 22, 4) {real, imag} */,
  {32'hc339e389, 32'hc2983d6e} /* (19, 22, 3) {real, imag} */,
  {32'h44797bab, 32'h42fe8bfa} /* (19, 22, 2) {real, imag} */,
  {32'hc511d2e7, 32'hc35b2428} /* (19, 22, 1) {real, imag} */,
  {32'hc525f4e9, 32'h00000000} /* (19, 22, 0) {real, imag} */,
  {32'hc43d92b0, 32'h42b9b040} /* (19, 21, 31) {real, imag} */,
  {32'h43d66136, 32'h421250e4} /* (19, 21, 30) {real, imag} */,
  {32'hc2aa6ff6, 32'h434a8d5c} /* (19, 21, 29) {real, imag} */,
  {32'hc2ddc98d, 32'hc2ee9b3b} /* (19, 21, 28) {real, imag} */,
  {32'h429e763c, 32'hc292740b} /* (19, 21, 27) {real, imag} */,
  {32'h4192396c, 32'h416b2a88} /* (19, 21, 26) {real, imag} */,
  {32'h41d76d46, 32'hc1fd2761} /* (19, 21, 25) {real, imag} */,
  {32'h424c8a08, 32'h41728196} /* (19, 21, 24) {real, imag} */,
  {32'h424a3cce, 32'h41c42464} /* (19, 21, 23) {real, imag} */,
  {32'hc1b9fd7a, 32'hc21ad586} /* (19, 21, 22) {real, imag} */,
  {32'hc11450a8, 32'h41c0f723} /* (19, 21, 21) {real, imag} */,
  {32'h41e3a296, 32'h42417c4a} /* (19, 21, 20) {real, imag} */,
  {32'hc1973a12, 32'hc0af2030} /* (19, 21, 19) {real, imag} */,
  {32'hc12ca214, 32'hc10b1740} /* (19, 21, 18) {real, imag} */,
  {32'h42483e96, 32'h401a0438} /* (19, 21, 17) {real, imag} */,
  {32'hc07c0390, 32'h00000000} /* (19, 21, 16) {real, imag} */,
  {32'h42483e96, 32'hc01a0438} /* (19, 21, 15) {real, imag} */,
  {32'hc12ca214, 32'h410b1740} /* (19, 21, 14) {real, imag} */,
  {32'hc1973a12, 32'h40af2030} /* (19, 21, 13) {real, imag} */,
  {32'h41e3a296, 32'hc2417c4a} /* (19, 21, 12) {real, imag} */,
  {32'hc11450a8, 32'hc1c0f723} /* (19, 21, 11) {real, imag} */,
  {32'hc1b9fd7a, 32'h421ad586} /* (19, 21, 10) {real, imag} */,
  {32'h424a3cce, 32'hc1c42464} /* (19, 21, 9) {real, imag} */,
  {32'h424c8a08, 32'hc1728196} /* (19, 21, 8) {real, imag} */,
  {32'h41d76d46, 32'h41fd2761} /* (19, 21, 7) {real, imag} */,
  {32'h4192396c, 32'hc16b2a88} /* (19, 21, 6) {real, imag} */,
  {32'h429e763c, 32'h4292740b} /* (19, 21, 5) {real, imag} */,
  {32'hc2ddc98d, 32'h42ee9b3b} /* (19, 21, 4) {real, imag} */,
  {32'hc2aa6ff6, 32'hc34a8d5c} /* (19, 21, 3) {real, imag} */,
  {32'h43d66136, 32'hc21250e4} /* (19, 21, 2) {real, imag} */,
  {32'hc43d92b0, 32'hc2b9b040} /* (19, 21, 1) {real, imag} */,
  {32'hc4a06f14, 32'h00000000} /* (19, 21, 0) {real, imag} */,
  {32'h448f4b07, 32'hc3729aa0} /* (19, 20, 31) {real, imag} */,
  {32'hc3c1062e, 32'h433cd662} /* (19, 20, 30) {real, imag} */,
  {32'hc2e93d46, 32'h421f8c6c} /* (19, 20, 29) {real, imag} */,
  {32'h43251ba0, 32'hc1892731} /* (19, 20, 28) {real, imag} */,
  {32'hc316bef8, 32'h430b13d5} /* (19, 20, 27) {real, imag} */,
  {32'h41f76758, 32'h42481cf9} /* (19, 20, 26) {real, imag} */,
  {32'h4302774e, 32'h4243db6a} /* (19, 20, 25) {real, imag} */,
  {32'hc2ca3a9d, 32'hc265e677} /* (19, 20, 24) {real, imag} */,
  {32'hc25f4bc4, 32'hc2d421bf} /* (19, 20, 23) {real, imag} */,
  {32'hc253653a, 32'hc1ad0c76} /* (19, 20, 22) {real, imag} */,
  {32'hc21466e4, 32'h4173b9d0} /* (19, 20, 21) {real, imag} */,
  {32'h42aa04f0, 32'hc1f1d622} /* (19, 20, 20) {real, imag} */,
  {32'h415dbf70, 32'h4276c852} /* (19, 20, 19) {real, imag} */,
  {32'hc004f1e8, 32'h42a19638} /* (19, 20, 18) {real, imag} */,
  {32'hc23f4a9d, 32'hc205a567} /* (19, 20, 17) {real, imag} */,
  {32'h42816546, 32'h00000000} /* (19, 20, 16) {real, imag} */,
  {32'hc23f4a9d, 32'h4205a567} /* (19, 20, 15) {real, imag} */,
  {32'hc004f1e8, 32'hc2a19638} /* (19, 20, 14) {real, imag} */,
  {32'h415dbf70, 32'hc276c852} /* (19, 20, 13) {real, imag} */,
  {32'h42aa04f0, 32'h41f1d622} /* (19, 20, 12) {real, imag} */,
  {32'hc21466e4, 32'hc173b9d0} /* (19, 20, 11) {real, imag} */,
  {32'hc253653a, 32'h41ad0c76} /* (19, 20, 10) {real, imag} */,
  {32'hc25f4bc4, 32'h42d421bf} /* (19, 20, 9) {real, imag} */,
  {32'hc2ca3a9d, 32'h4265e677} /* (19, 20, 8) {real, imag} */,
  {32'h4302774e, 32'hc243db6a} /* (19, 20, 7) {real, imag} */,
  {32'h41f76758, 32'hc2481cf9} /* (19, 20, 6) {real, imag} */,
  {32'hc316bef8, 32'hc30b13d5} /* (19, 20, 5) {real, imag} */,
  {32'h43251ba0, 32'h41892731} /* (19, 20, 4) {real, imag} */,
  {32'hc2e93d46, 32'hc21f8c6c} /* (19, 20, 3) {real, imag} */,
  {32'hc3c1062e, 32'hc33cd662} /* (19, 20, 2) {real, imag} */,
  {32'h448f4b07, 32'h43729aa0} /* (19, 20, 1) {real, imag} */,
  {32'h439412c0, 32'h00000000} /* (19, 20, 0) {real, imag} */,
  {32'h451cfe57, 32'hc3c45b00} /* (19, 19, 31) {real, imag} */,
  {32'hc469ca0c, 32'h42e798ba} /* (19, 19, 30) {real, imag} */,
  {32'hc1d4d7e6, 32'h431eeb1c} /* (19, 19, 29) {real, imag} */,
  {32'h437be862, 32'hc2604d63} /* (19, 19, 28) {real, imag} */,
  {32'hc3332efa, 32'h434bbe60} /* (19, 19, 27) {real, imag} */,
  {32'hc1cf52ea, 32'h42f62a7a} /* (19, 19, 26) {real, imag} */,
  {32'h4302f8ce, 32'hc26c96f2} /* (19, 19, 25) {real, imag} */,
  {32'h4260c6a8, 32'h42abf56c} /* (19, 19, 24) {real, imag} */,
  {32'h429da774, 32'hc2c90d06} /* (19, 19, 23) {real, imag} */,
  {32'hc2e2a386, 32'h4233a7f8} /* (19, 19, 22) {real, imag} */,
  {32'hc252d75a, 32'h4251c362} /* (19, 19, 21) {real, imag} */,
  {32'h4209d42e, 32'h4243e53a} /* (19, 19, 20) {real, imag} */,
  {32'hc22bf3cc, 32'hc22138ee} /* (19, 19, 19) {real, imag} */,
  {32'h40995698, 32'hc15acac0} /* (19, 19, 18) {real, imag} */,
  {32'h42649272, 32'h42417873} /* (19, 19, 17) {real, imag} */,
  {32'h42696b78, 32'h00000000} /* (19, 19, 16) {real, imag} */,
  {32'h42649272, 32'hc2417873} /* (19, 19, 15) {real, imag} */,
  {32'h40995698, 32'h415acac0} /* (19, 19, 14) {real, imag} */,
  {32'hc22bf3cc, 32'h422138ee} /* (19, 19, 13) {real, imag} */,
  {32'h4209d42e, 32'hc243e53a} /* (19, 19, 12) {real, imag} */,
  {32'hc252d75a, 32'hc251c362} /* (19, 19, 11) {real, imag} */,
  {32'hc2e2a386, 32'hc233a7f8} /* (19, 19, 10) {real, imag} */,
  {32'h429da774, 32'h42c90d06} /* (19, 19, 9) {real, imag} */,
  {32'h4260c6a8, 32'hc2abf56c} /* (19, 19, 8) {real, imag} */,
  {32'h4302f8ce, 32'h426c96f2} /* (19, 19, 7) {real, imag} */,
  {32'hc1cf52ea, 32'hc2f62a7a} /* (19, 19, 6) {real, imag} */,
  {32'hc3332efa, 32'hc34bbe60} /* (19, 19, 5) {real, imag} */,
  {32'h437be862, 32'h42604d63} /* (19, 19, 4) {real, imag} */,
  {32'hc1d4d7e6, 32'hc31eeb1c} /* (19, 19, 3) {real, imag} */,
  {32'hc469ca0c, 32'hc2e798ba} /* (19, 19, 2) {real, imag} */,
  {32'h451cfe57, 32'h43c45b00} /* (19, 19, 1) {real, imag} */,
  {32'h44b1175e, 32'h00000000} /* (19, 19, 0) {real, imag} */,
  {32'h45504838, 32'hc39bba90} /* (19, 18, 31) {real, imag} */,
  {32'hc4a3ee5e, 32'h43676b5b} /* (19, 18, 30) {real, imag} */,
  {32'h42fd5c78, 32'h4309bfd9} /* (19, 18, 29) {real, imag} */,
  {32'h439c2e78, 32'hc204da62} /* (19, 18, 28) {real, imag} */,
  {32'hc258d3ba, 32'h40f8c9f8} /* (19, 18, 27) {real, imag} */,
  {32'hc2aeec81, 32'hc32af88a} /* (19, 18, 26) {real, imag} */,
  {32'h4265ff0a, 32'h41b25188} /* (19, 18, 25) {real, imag} */,
  {32'h41cefc13, 32'h4311146f} /* (19, 18, 24) {real, imag} */,
  {32'h42e19d38, 32'hc2953670} /* (19, 18, 23) {real, imag} */,
  {32'h420d2e89, 32'h3f10a480} /* (19, 18, 22) {real, imag} */,
  {32'hc2e05188, 32'h431db0b0} /* (19, 18, 21) {real, imag} */,
  {32'hc1ad47a8, 32'h41ec1540} /* (19, 18, 20) {real, imag} */,
  {32'h42207679, 32'hc204a3eb} /* (19, 18, 19) {real, imag} */,
  {32'h42a03adc, 32'h423040bb} /* (19, 18, 18) {real, imag} */,
  {32'h4283c3b0, 32'h418dc00a} /* (19, 18, 17) {real, imag} */,
  {32'h408ca258, 32'h00000000} /* (19, 18, 16) {real, imag} */,
  {32'h4283c3b0, 32'hc18dc00a} /* (19, 18, 15) {real, imag} */,
  {32'h42a03adc, 32'hc23040bb} /* (19, 18, 14) {real, imag} */,
  {32'h42207679, 32'h4204a3eb} /* (19, 18, 13) {real, imag} */,
  {32'hc1ad47a8, 32'hc1ec1540} /* (19, 18, 12) {real, imag} */,
  {32'hc2e05188, 32'hc31db0b0} /* (19, 18, 11) {real, imag} */,
  {32'h420d2e89, 32'hbf10a480} /* (19, 18, 10) {real, imag} */,
  {32'h42e19d38, 32'h42953670} /* (19, 18, 9) {real, imag} */,
  {32'h41cefc13, 32'hc311146f} /* (19, 18, 8) {real, imag} */,
  {32'h4265ff0a, 32'hc1b25188} /* (19, 18, 7) {real, imag} */,
  {32'hc2aeec81, 32'h432af88a} /* (19, 18, 6) {real, imag} */,
  {32'hc258d3ba, 32'hc0f8c9f8} /* (19, 18, 5) {real, imag} */,
  {32'h439c2e78, 32'h4204da62} /* (19, 18, 4) {real, imag} */,
  {32'h42fd5c78, 32'hc309bfd9} /* (19, 18, 3) {real, imag} */,
  {32'hc4a3ee5e, 32'hc3676b5b} /* (19, 18, 2) {real, imag} */,
  {32'h45504838, 32'h439bba90} /* (19, 18, 1) {real, imag} */,
  {32'h4504e4a3, 32'h00000000} /* (19, 18, 0) {real, imag} */,
  {32'h456ca2ae, 32'hc3affe3f} /* (19, 17, 31) {real, imag} */,
  {32'hc4b7e339, 32'h437bf1ba} /* (19, 17, 30) {real, imag} */,
  {32'h41df7bba, 32'h42420f6a} /* (19, 17, 29) {real, imag} */,
  {32'h43149889, 32'hc2ba39ee} /* (19, 17, 28) {real, imag} */,
  {32'hc2b2203b, 32'h430f1aa4} /* (19, 17, 27) {real, imag} */,
  {32'hc2658b92, 32'hc02b7a50} /* (19, 17, 26) {real, imag} */,
  {32'h42f57412, 32'hc238691c} /* (19, 17, 25) {real, imag} */,
  {32'hc2c57b7d, 32'h42a282a8} /* (19, 17, 24) {real, imag} */,
  {32'h427c48ea, 32'h41aeb7c3} /* (19, 17, 23) {real, imag} */,
  {32'h3ead6ec0, 32'h42db3b6a} /* (19, 17, 22) {real, imag} */,
  {32'hc2050d64, 32'hc11a7995} /* (19, 17, 21) {real, imag} */,
  {32'h418a6c8e, 32'hc1c327aa} /* (19, 17, 20) {real, imag} */,
  {32'h42fb4665, 32'hc158f5b2} /* (19, 17, 19) {real, imag} */,
  {32'hc25ab622, 32'hc2ba4cf1} /* (19, 17, 18) {real, imag} */,
  {32'h4218e6db, 32'hc2c5c51a} /* (19, 17, 17) {real, imag} */,
  {32'h42b45098, 32'h00000000} /* (19, 17, 16) {real, imag} */,
  {32'h4218e6db, 32'h42c5c51a} /* (19, 17, 15) {real, imag} */,
  {32'hc25ab622, 32'h42ba4cf1} /* (19, 17, 14) {real, imag} */,
  {32'h42fb4665, 32'h4158f5b2} /* (19, 17, 13) {real, imag} */,
  {32'h418a6c8e, 32'h41c327aa} /* (19, 17, 12) {real, imag} */,
  {32'hc2050d64, 32'h411a7995} /* (19, 17, 11) {real, imag} */,
  {32'h3ead6ec0, 32'hc2db3b6a} /* (19, 17, 10) {real, imag} */,
  {32'h427c48ea, 32'hc1aeb7c3} /* (19, 17, 9) {real, imag} */,
  {32'hc2c57b7d, 32'hc2a282a8} /* (19, 17, 8) {real, imag} */,
  {32'h42f57412, 32'h4238691c} /* (19, 17, 7) {real, imag} */,
  {32'hc2658b92, 32'h402b7a50} /* (19, 17, 6) {real, imag} */,
  {32'hc2b2203b, 32'hc30f1aa4} /* (19, 17, 5) {real, imag} */,
  {32'h43149889, 32'h42ba39ee} /* (19, 17, 4) {real, imag} */,
  {32'h41df7bba, 32'hc2420f6a} /* (19, 17, 3) {real, imag} */,
  {32'hc4b7e339, 32'hc37bf1ba} /* (19, 17, 2) {real, imag} */,
  {32'h456ca2ae, 32'h43affe3f} /* (19, 17, 1) {real, imag} */,
  {32'h45276c76, 32'h00000000} /* (19, 17, 0) {real, imag} */,
  {32'h457c2b48, 32'hc3c1394c} /* (19, 16, 31) {real, imag} */,
  {32'hc4d00f64, 32'h4304b824} /* (19, 16, 30) {real, imag} */,
  {32'hc2c29584, 32'hc1b466b5} /* (19, 16, 29) {real, imag} */,
  {32'h438875dc, 32'hc21ac301} /* (19, 16, 28) {real, imag} */,
  {32'hc3458731, 32'h4314bd42} /* (19, 16, 27) {real, imag} */,
  {32'hc2924f74, 32'h4192180f} /* (19, 16, 26) {real, imag} */,
  {32'h4222465f, 32'hc2859075} /* (19, 16, 25) {real, imag} */,
  {32'hc227b5d9, 32'h41f75a2b} /* (19, 16, 24) {real, imag} */,
  {32'hc137cc54, 32'hc2c01b18} /* (19, 16, 23) {real, imag} */,
  {32'h3f99885c, 32'hc2d93e24} /* (19, 16, 22) {real, imag} */,
  {32'hc2982e39, 32'h42cf2077} /* (19, 16, 21) {real, imag} */,
  {32'hc225deb6, 32'h41e91206} /* (19, 16, 20) {real, imag} */,
  {32'hc2278c9d, 32'hc2d05555} /* (19, 16, 19) {real, imag} */,
  {32'h40821344, 32'h4259e2c2} /* (19, 16, 18) {real, imag} */,
  {32'hc27cd8e6, 32'hc233e872} /* (19, 16, 17) {real, imag} */,
  {32'hc1efffbc, 32'h00000000} /* (19, 16, 16) {real, imag} */,
  {32'hc27cd8e6, 32'h4233e872} /* (19, 16, 15) {real, imag} */,
  {32'h40821344, 32'hc259e2c2} /* (19, 16, 14) {real, imag} */,
  {32'hc2278c9d, 32'h42d05555} /* (19, 16, 13) {real, imag} */,
  {32'hc225deb6, 32'hc1e91206} /* (19, 16, 12) {real, imag} */,
  {32'hc2982e39, 32'hc2cf2077} /* (19, 16, 11) {real, imag} */,
  {32'h3f99885c, 32'h42d93e24} /* (19, 16, 10) {real, imag} */,
  {32'hc137cc54, 32'h42c01b18} /* (19, 16, 9) {real, imag} */,
  {32'hc227b5d9, 32'hc1f75a2b} /* (19, 16, 8) {real, imag} */,
  {32'h4222465f, 32'h42859075} /* (19, 16, 7) {real, imag} */,
  {32'hc2924f74, 32'hc192180f} /* (19, 16, 6) {real, imag} */,
  {32'hc3458731, 32'hc314bd42} /* (19, 16, 5) {real, imag} */,
  {32'h438875dc, 32'h421ac301} /* (19, 16, 4) {real, imag} */,
  {32'hc2c29584, 32'h41b466b5} /* (19, 16, 3) {real, imag} */,
  {32'hc4d00f64, 32'hc304b824} /* (19, 16, 2) {real, imag} */,
  {32'h457c2b48, 32'h43c1394c} /* (19, 16, 1) {real, imag} */,
  {32'h452e858c, 32'h00000000} /* (19, 16, 0) {real, imag} */,
  {32'h457b1aee, 32'hc3b54321} /* (19, 15, 31) {real, imag} */,
  {32'hc4e08491, 32'h435f4d46} /* (19, 15, 30) {real, imag} */,
  {32'hc2230f1f, 32'hc2486828} /* (19, 15, 29) {real, imag} */,
  {32'h43b3a454, 32'hc2cf0cd2} /* (19, 15, 28) {real, imag} */,
  {32'hc355ca22, 32'h430c1d30} /* (19, 15, 27) {real, imag} */,
  {32'hc19b31a4, 32'h4135210c} /* (19, 15, 26) {real, imag} */,
  {32'hc1de1a66, 32'hc2f2d27a} /* (19, 15, 25) {real, imag} */,
  {32'h416b46c8, 32'h42ad4c4a} /* (19, 15, 24) {real, imag} */,
  {32'hc297631d, 32'hc202ec9e} /* (19, 15, 23) {real, imag} */,
  {32'h3fb0f370, 32'h4205e8cb} /* (19, 15, 22) {real, imag} */,
  {32'hc1a6c347, 32'h4224fbc7} /* (19, 15, 21) {real, imag} */,
  {32'hc2a1cc52, 32'hc291febc} /* (19, 15, 20) {real, imag} */,
  {32'h41227b38, 32'h41a65ae7} /* (19, 15, 19) {real, imag} */,
  {32'hc121f1c6, 32'h42fb285b} /* (19, 15, 18) {real, imag} */,
  {32'hc22db9b7, 32'h4065b2c0} /* (19, 15, 17) {real, imag} */,
  {32'h42bfd88a, 32'h00000000} /* (19, 15, 16) {real, imag} */,
  {32'hc22db9b7, 32'hc065b2c0} /* (19, 15, 15) {real, imag} */,
  {32'hc121f1c6, 32'hc2fb285b} /* (19, 15, 14) {real, imag} */,
  {32'h41227b38, 32'hc1a65ae7} /* (19, 15, 13) {real, imag} */,
  {32'hc2a1cc52, 32'h4291febc} /* (19, 15, 12) {real, imag} */,
  {32'hc1a6c347, 32'hc224fbc7} /* (19, 15, 11) {real, imag} */,
  {32'h3fb0f370, 32'hc205e8cb} /* (19, 15, 10) {real, imag} */,
  {32'hc297631d, 32'h4202ec9e} /* (19, 15, 9) {real, imag} */,
  {32'h416b46c8, 32'hc2ad4c4a} /* (19, 15, 8) {real, imag} */,
  {32'hc1de1a66, 32'h42f2d27a} /* (19, 15, 7) {real, imag} */,
  {32'hc19b31a4, 32'hc135210c} /* (19, 15, 6) {real, imag} */,
  {32'hc355ca22, 32'hc30c1d30} /* (19, 15, 5) {real, imag} */,
  {32'h43b3a454, 32'h42cf0cd2} /* (19, 15, 4) {real, imag} */,
  {32'hc2230f1f, 32'h42486828} /* (19, 15, 3) {real, imag} */,
  {32'hc4e08491, 32'hc35f4d46} /* (19, 15, 2) {real, imag} */,
  {32'h457b1aee, 32'h43b54321} /* (19, 15, 1) {real, imag} */,
  {32'h453c209e, 32'h00000000} /* (19, 15, 0) {real, imag} */,
  {32'h4565f46a, 32'hc39335f0} /* (19, 14, 31) {real, imag} */,
  {32'hc4cf520a, 32'h4379245d} /* (19, 14, 30) {real, imag} */,
  {32'h422ab667, 32'hc1b98980} /* (19, 14, 29) {real, imag} */,
  {32'h432815f9, 32'hc295e927} /* (19, 14, 28) {real, imag} */,
  {32'hc35fb7e6, 32'h42aa9b6c} /* (19, 14, 27) {real, imag} */,
  {32'hc2a13975, 32'h430ad832} /* (19, 14, 26) {real, imag} */,
  {32'h421e9cea, 32'hc2c5e585} /* (19, 14, 25) {real, imag} */,
  {32'hc13e259e, 32'h42c06c7f} /* (19, 14, 24) {real, imag} */,
  {32'h42899b94, 32'hc2317fba} /* (19, 14, 23) {real, imag} */,
  {32'hc227b1d5, 32'hc29e6667} /* (19, 14, 22) {real, imag} */,
  {32'hc1d34832, 32'h424b4558} /* (19, 14, 21) {real, imag} */,
  {32'hbf2622c0, 32'h413dfd60} /* (19, 14, 20) {real, imag} */,
  {32'hc204777f, 32'h41c7ac78} /* (19, 14, 19) {real, imag} */,
  {32'hc264c0f8, 32'hc05daf20} /* (19, 14, 18) {real, imag} */,
  {32'h41929348, 32'h4221346d} /* (19, 14, 17) {real, imag} */,
  {32'h425c0185, 32'h00000000} /* (19, 14, 16) {real, imag} */,
  {32'h41929348, 32'hc221346d} /* (19, 14, 15) {real, imag} */,
  {32'hc264c0f8, 32'h405daf20} /* (19, 14, 14) {real, imag} */,
  {32'hc204777f, 32'hc1c7ac78} /* (19, 14, 13) {real, imag} */,
  {32'hbf2622c0, 32'hc13dfd60} /* (19, 14, 12) {real, imag} */,
  {32'hc1d34832, 32'hc24b4558} /* (19, 14, 11) {real, imag} */,
  {32'hc227b1d5, 32'h429e6667} /* (19, 14, 10) {real, imag} */,
  {32'h42899b94, 32'h42317fba} /* (19, 14, 9) {real, imag} */,
  {32'hc13e259e, 32'hc2c06c7f} /* (19, 14, 8) {real, imag} */,
  {32'h421e9cea, 32'h42c5e585} /* (19, 14, 7) {real, imag} */,
  {32'hc2a13975, 32'hc30ad832} /* (19, 14, 6) {real, imag} */,
  {32'hc35fb7e6, 32'hc2aa9b6c} /* (19, 14, 5) {real, imag} */,
  {32'h432815f9, 32'h4295e927} /* (19, 14, 4) {real, imag} */,
  {32'h422ab667, 32'h41b98980} /* (19, 14, 3) {real, imag} */,
  {32'hc4cf520a, 32'hc379245d} /* (19, 14, 2) {real, imag} */,
  {32'h4565f46a, 32'h439335f0} /* (19, 14, 1) {real, imag} */,
  {32'h452490b1, 32'h00000000} /* (19, 14, 0) {real, imag} */,
  {32'h4541aae5, 32'hc2fdf460} /* (19, 13, 31) {real, imag} */,
  {32'hc4b21a66, 32'h4345fc9f} /* (19, 13, 30) {real, imag} */,
  {32'h4282ccb0, 32'hc377321c} /* (19, 13, 29) {real, imag} */,
  {32'h43235e2e, 32'hc1d5f32a} /* (19, 13, 28) {real, imag} */,
  {32'hc36ca15e, 32'h41ba5020} /* (19, 13, 27) {real, imag} */,
  {32'h42536827, 32'h42a9e68e} /* (19, 13, 26) {real, imag} */,
  {32'hc23fe7d2, 32'hc1ec28d4} /* (19, 13, 25) {real, imag} */,
  {32'hc1e68118, 32'h420bb74c} /* (19, 13, 24) {real, imag} */,
  {32'h429796f0, 32'h41baa050} /* (19, 13, 23) {real, imag} */,
  {32'hc2ae5e3e, 32'hc302e785} /* (19, 13, 22) {real, imag} */,
  {32'hc21fa3cc, 32'h42a55cdb} /* (19, 13, 21) {real, imag} */,
  {32'h421fac28, 32'hc1d3286d} /* (19, 13, 20) {real, imag} */,
  {32'hc1d5135c, 32'h418e52d1} /* (19, 13, 19) {real, imag} */,
  {32'h42c4c888, 32'h4313cb53} /* (19, 13, 18) {real, imag} */,
  {32'h41e6bd04, 32'hc22a30c3} /* (19, 13, 17) {real, imag} */,
  {32'h42856cec, 32'h00000000} /* (19, 13, 16) {real, imag} */,
  {32'h41e6bd04, 32'h422a30c3} /* (19, 13, 15) {real, imag} */,
  {32'h42c4c888, 32'hc313cb53} /* (19, 13, 14) {real, imag} */,
  {32'hc1d5135c, 32'hc18e52d1} /* (19, 13, 13) {real, imag} */,
  {32'h421fac28, 32'h41d3286d} /* (19, 13, 12) {real, imag} */,
  {32'hc21fa3cc, 32'hc2a55cdb} /* (19, 13, 11) {real, imag} */,
  {32'hc2ae5e3e, 32'h4302e785} /* (19, 13, 10) {real, imag} */,
  {32'h429796f0, 32'hc1baa050} /* (19, 13, 9) {real, imag} */,
  {32'hc1e68118, 32'hc20bb74c} /* (19, 13, 8) {real, imag} */,
  {32'hc23fe7d2, 32'h41ec28d4} /* (19, 13, 7) {real, imag} */,
  {32'h42536827, 32'hc2a9e68e} /* (19, 13, 6) {real, imag} */,
  {32'hc36ca15e, 32'hc1ba5020} /* (19, 13, 5) {real, imag} */,
  {32'h43235e2e, 32'h41d5f32a} /* (19, 13, 4) {real, imag} */,
  {32'h4282ccb0, 32'h4377321c} /* (19, 13, 3) {real, imag} */,
  {32'hc4b21a66, 32'hc345fc9f} /* (19, 13, 2) {real, imag} */,
  {32'h4541aae5, 32'h42fdf460} /* (19, 13, 1) {real, imag} */,
  {32'h4503b053, 32'h00000000} /* (19, 13, 0) {real, imag} */,
  {32'h45082968, 32'h4270a980} /* (19, 12, 31) {real, imag} */,
  {32'hc49bb6e6, 32'h4387dfa8} /* (19, 12, 30) {real, imag} */,
  {32'h43158b45, 32'hc34019d1} /* (19, 12, 29) {real, imag} */,
  {32'h42c32859, 32'hc1bd6071} /* (19, 12, 28) {real, imag} */,
  {32'hc3625364, 32'h4324f16f} /* (19, 12, 27) {real, imag} */,
  {32'h42beafca, 32'h421b378f} /* (19, 12, 26) {real, imag} */,
  {32'hc23f2fca, 32'hc1e2357c} /* (19, 12, 25) {real, imag} */,
  {32'hc2ef7953, 32'hc1c53582} /* (19, 12, 24) {real, imag} */,
  {32'h419b9f58, 32'h42f05f21} /* (19, 12, 23) {real, imag} */,
  {32'hbf037e00, 32'hc244e217} /* (19, 12, 22) {real, imag} */,
  {32'h41f64c3f, 32'h420cafb8} /* (19, 12, 21) {real, imag} */,
  {32'h423ead11, 32'hc27e420d} /* (19, 12, 20) {real, imag} */,
  {32'hc2733ea0, 32'h42b77431} /* (19, 12, 19) {real, imag} */,
  {32'h42728f94, 32'h41d02c38} /* (19, 12, 18) {real, imag} */,
  {32'hc2238cb9, 32'hc15f9f80} /* (19, 12, 17) {real, imag} */,
  {32'hc1b7d42a, 32'h00000000} /* (19, 12, 16) {real, imag} */,
  {32'hc2238cb9, 32'h415f9f80} /* (19, 12, 15) {real, imag} */,
  {32'h42728f94, 32'hc1d02c38} /* (19, 12, 14) {real, imag} */,
  {32'hc2733ea0, 32'hc2b77431} /* (19, 12, 13) {real, imag} */,
  {32'h423ead11, 32'h427e420d} /* (19, 12, 12) {real, imag} */,
  {32'h41f64c3f, 32'hc20cafb8} /* (19, 12, 11) {real, imag} */,
  {32'hbf037e00, 32'h4244e217} /* (19, 12, 10) {real, imag} */,
  {32'h419b9f58, 32'hc2f05f21} /* (19, 12, 9) {real, imag} */,
  {32'hc2ef7953, 32'h41c53582} /* (19, 12, 8) {real, imag} */,
  {32'hc23f2fca, 32'h41e2357c} /* (19, 12, 7) {real, imag} */,
  {32'h42beafca, 32'hc21b378f} /* (19, 12, 6) {real, imag} */,
  {32'hc3625364, 32'hc324f16f} /* (19, 12, 5) {real, imag} */,
  {32'h42c32859, 32'h41bd6071} /* (19, 12, 4) {real, imag} */,
  {32'h43158b45, 32'h434019d1} /* (19, 12, 3) {real, imag} */,
  {32'hc49bb6e6, 32'hc387dfa8} /* (19, 12, 2) {real, imag} */,
  {32'h45082968, 32'hc270a980} /* (19, 12, 1) {real, imag} */,
  {32'h44b3c06e, 32'h00000000} /* (19, 12, 0) {real, imag} */,
  {32'h44736eb0, 32'h43abbdf8} /* (19, 11, 31) {real, imag} */,
  {32'hc41b3e2d, 32'h42c59906} /* (19, 11, 30) {real, imag} */,
  {32'h430608c8, 32'hc2b52d08} /* (19, 11, 29) {real, imag} */,
  {32'h42c2e0a3, 32'hc0f425a0} /* (19, 11, 28) {real, imag} */,
  {32'hc3722a6e, 32'h41a44704} /* (19, 11, 27) {real, imag} */,
  {32'h42f1e0d9, 32'h418d5ac8} /* (19, 11, 26) {real, imag} */,
  {32'hc2ec53ae, 32'h4226eb76} /* (19, 11, 25) {real, imag} */,
  {32'hc296422f, 32'hc1d29903} /* (19, 11, 24) {real, imag} */,
  {32'h4239dee0, 32'h4207dcfa} /* (19, 11, 23) {real, imag} */,
  {32'hc105b91c, 32'hc2a68399} /* (19, 11, 22) {real, imag} */,
  {32'hc2719c58, 32'h416573ba} /* (19, 11, 21) {real, imag} */,
  {32'h42904d70, 32'h404bb7c8} /* (19, 11, 20) {real, imag} */,
  {32'hc05baef4, 32'h42a7b567} /* (19, 11, 19) {real, imag} */,
  {32'h41dfc734, 32'hc1ae8a78} /* (19, 11, 18) {real, imag} */,
  {32'h409ed9fc, 32'h425185aa} /* (19, 11, 17) {real, imag} */,
  {32'h42d4dbc8, 32'h00000000} /* (19, 11, 16) {real, imag} */,
  {32'h409ed9fc, 32'hc25185aa} /* (19, 11, 15) {real, imag} */,
  {32'h41dfc734, 32'h41ae8a78} /* (19, 11, 14) {real, imag} */,
  {32'hc05baef4, 32'hc2a7b567} /* (19, 11, 13) {real, imag} */,
  {32'h42904d70, 32'hc04bb7c8} /* (19, 11, 12) {real, imag} */,
  {32'hc2719c58, 32'hc16573ba} /* (19, 11, 11) {real, imag} */,
  {32'hc105b91c, 32'h42a68399} /* (19, 11, 10) {real, imag} */,
  {32'h4239dee0, 32'hc207dcfa} /* (19, 11, 9) {real, imag} */,
  {32'hc296422f, 32'h41d29903} /* (19, 11, 8) {real, imag} */,
  {32'hc2ec53ae, 32'hc226eb76} /* (19, 11, 7) {real, imag} */,
  {32'h42f1e0d9, 32'hc18d5ac8} /* (19, 11, 6) {real, imag} */,
  {32'hc3722a6e, 32'hc1a44704} /* (19, 11, 5) {real, imag} */,
  {32'h42c2e0a3, 32'h40f425a0} /* (19, 11, 4) {real, imag} */,
  {32'h430608c8, 32'h42b52d08} /* (19, 11, 3) {real, imag} */,
  {32'hc41b3e2d, 32'hc2c59906} /* (19, 11, 2) {real, imag} */,
  {32'h44736eb0, 32'hc3abbdf8} /* (19, 11, 1) {real, imag} */,
  {32'h44088258, 32'h00000000} /* (19, 11, 0) {real, imag} */,
  {32'hc45cbab1, 32'h44490ab8} /* (19, 10, 31) {real, imag} */,
  {32'h43b8218a, 32'hc2af0352} /* (19, 10, 30) {real, imag} */,
  {32'hbf5bcd00, 32'hc29e78b2} /* (19, 10, 29) {real, imag} */,
  {32'hc27cccbe, 32'h40628e30} /* (19, 10, 28) {real, imag} */,
  {32'hc0819bc0, 32'h41a74d30} /* (19, 10, 27) {real, imag} */,
  {32'h429bcd3a, 32'hc25bd378} /* (19, 10, 26) {real, imag} */,
  {32'hc3056f96, 32'h42d27b2c} /* (19, 10, 25) {real, imag} */,
  {32'hc1369ffc, 32'hc2c31244} /* (19, 10, 24) {real, imag} */,
  {32'h424c59ac, 32'h430ef52b} /* (19, 10, 23) {real, imag} */,
  {32'h42873efc, 32'hc17a2752} /* (19, 10, 22) {real, imag} */,
  {32'hc1ac60b4, 32'h42606766} /* (19, 10, 21) {real, imag} */,
  {32'hc21bffe4, 32'hc125dcac} /* (19, 10, 20) {real, imag} */,
  {32'h41e0d77e, 32'hc18a373b} /* (19, 10, 19) {real, imag} */,
  {32'h41bbd08c, 32'h4206c71a} /* (19, 10, 18) {real, imag} */,
  {32'hc1e5141f, 32'hc29bf14e} /* (19, 10, 17) {real, imag} */,
  {32'h4221c48c, 32'h00000000} /* (19, 10, 16) {real, imag} */,
  {32'hc1e5141f, 32'h429bf14e} /* (19, 10, 15) {real, imag} */,
  {32'h41bbd08c, 32'hc206c71a} /* (19, 10, 14) {real, imag} */,
  {32'h41e0d77e, 32'h418a373b} /* (19, 10, 13) {real, imag} */,
  {32'hc21bffe4, 32'h4125dcac} /* (19, 10, 12) {real, imag} */,
  {32'hc1ac60b4, 32'hc2606766} /* (19, 10, 11) {real, imag} */,
  {32'h42873efc, 32'h417a2752} /* (19, 10, 10) {real, imag} */,
  {32'h424c59ac, 32'hc30ef52b} /* (19, 10, 9) {real, imag} */,
  {32'hc1369ffc, 32'h42c31244} /* (19, 10, 8) {real, imag} */,
  {32'hc3056f96, 32'hc2d27b2c} /* (19, 10, 7) {real, imag} */,
  {32'h429bcd3a, 32'h425bd378} /* (19, 10, 6) {real, imag} */,
  {32'hc0819bc0, 32'hc1a74d30} /* (19, 10, 5) {real, imag} */,
  {32'hc27cccbe, 32'hc0628e30} /* (19, 10, 4) {real, imag} */,
  {32'hbf5bcd00, 32'h429e78b2} /* (19, 10, 3) {real, imag} */,
  {32'h43b8218a, 32'h42af0352} /* (19, 10, 2) {real, imag} */,
  {32'hc45cbab1, 32'hc4490ab8} /* (19, 10, 1) {real, imag} */,
  {32'hc462157c, 32'h00000000} /* (19, 10, 0) {real, imag} */,
  {32'hc51164b1, 32'h44840e23} /* (19, 9, 31) {real, imag} */,
  {32'h446db53c, 32'hc356dd12} /* (19, 9, 30) {real, imag} */,
  {32'hc30b43ca, 32'h41c786b8} /* (19, 9, 29) {real, imag} */,
  {32'h41e99f74, 32'hc1d0d088} /* (19, 9, 28) {real, imag} */,
  {32'h42c3ca6a, 32'h4189f190} /* (19, 9, 27) {real, imag} */,
  {32'h41c50728, 32'hc249743a} /* (19, 9, 26) {real, imag} */,
  {32'hc33a21e9, 32'h420727c0} /* (19, 9, 25) {real, imag} */,
  {32'h426a6f40, 32'hc30f0faf} /* (19, 9, 24) {real, imag} */,
  {32'h428002ab, 32'h42a15320} /* (19, 9, 23) {real, imag} */,
  {32'hc304238a, 32'h41e7bfb0} /* (19, 9, 22) {real, imag} */,
  {32'h42d42a09, 32'hc2631a3c} /* (19, 9, 21) {real, imag} */,
  {32'hc002c2a4, 32'hc218caea} /* (19, 9, 20) {real, imag} */,
  {32'h43294946, 32'hc24f2d3d} /* (19, 9, 19) {real, imag} */,
  {32'hc3010c1f, 32'hc20717cb} /* (19, 9, 18) {real, imag} */,
  {32'hc2418624, 32'hc11ecc42} /* (19, 9, 17) {real, imag} */,
  {32'hc2611c59, 32'h00000000} /* (19, 9, 16) {real, imag} */,
  {32'hc2418624, 32'h411ecc42} /* (19, 9, 15) {real, imag} */,
  {32'hc3010c1f, 32'h420717cb} /* (19, 9, 14) {real, imag} */,
  {32'h43294946, 32'h424f2d3d} /* (19, 9, 13) {real, imag} */,
  {32'hc002c2a4, 32'h4218caea} /* (19, 9, 12) {real, imag} */,
  {32'h42d42a09, 32'h42631a3c} /* (19, 9, 11) {real, imag} */,
  {32'hc304238a, 32'hc1e7bfb0} /* (19, 9, 10) {real, imag} */,
  {32'h428002ab, 32'hc2a15320} /* (19, 9, 9) {real, imag} */,
  {32'h426a6f40, 32'h430f0faf} /* (19, 9, 8) {real, imag} */,
  {32'hc33a21e9, 32'hc20727c0} /* (19, 9, 7) {real, imag} */,
  {32'h41c50728, 32'h4249743a} /* (19, 9, 6) {real, imag} */,
  {32'h42c3ca6a, 32'hc189f190} /* (19, 9, 5) {real, imag} */,
  {32'h41e99f74, 32'h41d0d088} /* (19, 9, 4) {real, imag} */,
  {32'hc30b43ca, 32'hc1c786b8} /* (19, 9, 3) {real, imag} */,
  {32'h446db53c, 32'h4356dd12} /* (19, 9, 2) {real, imag} */,
  {32'hc51164b1, 32'hc4840e23} /* (19, 9, 1) {real, imag} */,
  {32'hc4f7d4a4, 32'h00000000} /* (19, 9, 0) {real, imag} */,
  {32'hc53ffaa7, 32'h44ad88fb} /* (19, 8, 31) {real, imag} */,
  {32'h4476cc3e, 32'hc3912a5c} /* (19, 8, 30) {real, imag} */,
  {32'hc2b411c1, 32'hc01b04d8} /* (19, 8, 29) {real, imag} */,
  {32'hc2f76aa6, 32'h4225af66} /* (19, 8, 28) {real, imag} */,
  {32'h4344ff42, 32'hc2307d97} /* (19, 8, 27) {real, imag} */,
  {32'hc242e0e9, 32'hc278e0ee} /* (19, 8, 26) {real, imag} */,
  {32'hc21f416a, 32'h41518978} /* (19, 8, 25) {real, imag} */,
  {32'h42cfe75a, 32'hc2865aea} /* (19, 8, 24) {real, imag} */,
  {32'h429bb450, 32'h429ed10a} /* (19, 8, 23) {real, imag} */,
  {32'hc32bb4ff, 32'hc1b3ad39} /* (19, 8, 22) {real, imag} */,
  {32'hc1508450, 32'hc32fe75e} /* (19, 8, 21) {real, imag} */,
  {32'hc232c308, 32'hc11e033a} /* (19, 8, 20) {real, imag} */,
  {32'hc2068084, 32'h41a38cee} /* (19, 8, 19) {real, imag} */,
  {32'h4175fb76, 32'hc2833a9a} /* (19, 8, 18) {real, imag} */,
  {32'h4279782b, 32'h4183a83c} /* (19, 8, 17) {real, imag} */,
  {32'hc137dc90, 32'h00000000} /* (19, 8, 16) {real, imag} */,
  {32'h4279782b, 32'hc183a83c} /* (19, 8, 15) {real, imag} */,
  {32'h4175fb76, 32'h42833a9a} /* (19, 8, 14) {real, imag} */,
  {32'hc2068084, 32'hc1a38cee} /* (19, 8, 13) {real, imag} */,
  {32'hc232c308, 32'h411e033a} /* (19, 8, 12) {real, imag} */,
  {32'hc1508450, 32'h432fe75e} /* (19, 8, 11) {real, imag} */,
  {32'hc32bb4ff, 32'h41b3ad39} /* (19, 8, 10) {real, imag} */,
  {32'h429bb450, 32'hc29ed10a} /* (19, 8, 9) {real, imag} */,
  {32'h42cfe75a, 32'h42865aea} /* (19, 8, 8) {real, imag} */,
  {32'hc21f416a, 32'hc1518978} /* (19, 8, 7) {real, imag} */,
  {32'hc242e0e9, 32'h4278e0ee} /* (19, 8, 6) {real, imag} */,
  {32'h4344ff42, 32'h42307d97} /* (19, 8, 5) {real, imag} */,
  {32'hc2f76aa6, 32'hc225af66} /* (19, 8, 4) {real, imag} */,
  {32'hc2b411c1, 32'h401b04d8} /* (19, 8, 3) {real, imag} */,
  {32'h4476cc3e, 32'h43912a5c} /* (19, 8, 2) {real, imag} */,
  {32'hc53ffaa7, 32'hc4ad88fb} /* (19, 8, 1) {real, imag} */,
  {32'hc533073c, 32'h00000000} /* (19, 8, 0) {real, imag} */,
  {32'hc559fd84, 32'h44e874ee} /* (19, 7, 31) {real, imag} */,
  {32'h44861c1c, 32'hc406d418} /* (19, 7, 30) {real, imag} */,
  {32'hc30a43d3, 32'hc08c1de8} /* (19, 7, 29) {real, imag} */,
  {32'hc2ca1cc0, 32'h431b6b27} /* (19, 7, 28) {real, imag} */,
  {32'h430929a3, 32'hc25be488} /* (19, 7, 27) {real, imag} */,
  {32'hc15fe1a4, 32'h422eea88} /* (19, 7, 26) {real, imag} */,
  {32'h42a84f6c, 32'h42787926} /* (19, 7, 25) {real, imag} */,
  {32'hc197bc12, 32'hc2f892d6} /* (19, 7, 24) {real, imag} */,
  {32'hc204f7ce, 32'h42ca3106} /* (19, 7, 23) {real, imag} */,
  {32'h428537e4, 32'h4292a014} /* (19, 7, 22) {real, imag} */,
  {32'h42ea81da, 32'hc3015eec} /* (19, 7, 21) {real, imag} */,
  {32'hc26b0066, 32'h42be7140} /* (19, 7, 20) {real, imag} */,
  {32'hc0b8a970, 32'h42ca7637} /* (19, 7, 19) {real, imag} */,
  {32'h41588c96, 32'h419e8e48} /* (19, 7, 18) {real, imag} */,
  {32'h420f3f9a, 32'h421a0a8c} /* (19, 7, 17) {real, imag} */,
  {32'hc23385dc, 32'h00000000} /* (19, 7, 16) {real, imag} */,
  {32'h420f3f9a, 32'hc21a0a8c} /* (19, 7, 15) {real, imag} */,
  {32'h41588c96, 32'hc19e8e48} /* (19, 7, 14) {real, imag} */,
  {32'hc0b8a970, 32'hc2ca7637} /* (19, 7, 13) {real, imag} */,
  {32'hc26b0066, 32'hc2be7140} /* (19, 7, 12) {real, imag} */,
  {32'h42ea81da, 32'h43015eec} /* (19, 7, 11) {real, imag} */,
  {32'h428537e4, 32'hc292a014} /* (19, 7, 10) {real, imag} */,
  {32'hc204f7ce, 32'hc2ca3106} /* (19, 7, 9) {real, imag} */,
  {32'hc197bc12, 32'h42f892d6} /* (19, 7, 8) {real, imag} */,
  {32'h42a84f6c, 32'hc2787926} /* (19, 7, 7) {real, imag} */,
  {32'hc15fe1a4, 32'hc22eea88} /* (19, 7, 6) {real, imag} */,
  {32'h430929a3, 32'h425be488} /* (19, 7, 5) {real, imag} */,
  {32'hc2ca1cc0, 32'hc31b6b27} /* (19, 7, 4) {real, imag} */,
  {32'hc30a43d3, 32'h408c1de8} /* (19, 7, 3) {real, imag} */,
  {32'h44861c1c, 32'h4406d418} /* (19, 7, 2) {real, imag} */,
  {32'hc559fd84, 32'hc4e874ee} /* (19, 7, 1) {real, imag} */,
  {32'hc560e3ce, 32'h00000000} /* (19, 7, 0) {real, imag} */,
  {32'hc56123f8, 32'h4507f18b} /* (19, 6, 31) {real, imag} */,
  {32'h44538b6f, 32'hc438faac} /* (19, 6, 30) {real, imag} */,
  {32'hc2922014, 32'hc2819ca5} /* (19, 6, 29) {real, imag} */,
  {32'hc2281bc0, 32'hbdedc200} /* (19, 6, 28) {real, imag} */,
  {32'h42deb268, 32'hc19e10b0} /* (19, 6, 27) {real, imag} */,
  {32'h3fc7c980, 32'h4115bf18} /* (19, 6, 26) {real, imag} */,
  {32'h4318d48a, 32'hc194ddea} /* (19, 6, 25) {real, imag} */,
  {32'h41acc0fc, 32'hc32c5aa2} /* (19, 6, 24) {real, imag} */,
  {32'hc0fe3cfa, 32'hc226520e} /* (19, 6, 23) {real, imag} */,
  {32'hc25f4c48, 32'h42cb4f03} /* (19, 6, 22) {real, imag} */,
  {32'h415eddb8, 32'hc1e0a6c8} /* (19, 6, 21) {real, imag} */,
  {32'hc27631e1, 32'h411ed667} /* (19, 6, 20) {real, imag} */,
  {32'h42456a70, 32'hc24ead7c} /* (19, 6, 19) {real, imag} */,
  {32'h430105b0, 32'hc21793fa} /* (19, 6, 18) {real, imag} */,
  {32'hc25eda06, 32'hc09882ba} /* (19, 6, 17) {real, imag} */,
  {32'h411efe0f, 32'h00000000} /* (19, 6, 16) {real, imag} */,
  {32'hc25eda06, 32'h409882ba} /* (19, 6, 15) {real, imag} */,
  {32'h430105b0, 32'h421793fa} /* (19, 6, 14) {real, imag} */,
  {32'h42456a70, 32'h424ead7c} /* (19, 6, 13) {real, imag} */,
  {32'hc27631e1, 32'hc11ed667} /* (19, 6, 12) {real, imag} */,
  {32'h415eddb8, 32'h41e0a6c8} /* (19, 6, 11) {real, imag} */,
  {32'hc25f4c48, 32'hc2cb4f03} /* (19, 6, 10) {real, imag} */,
  {32'hc0fe3cfa, 32'h4226520e} /* (19, 6, 9) {real, imag} */,
  {32'h41acc0fc, 32'h432c5aa2} /* (19, 6, 8) {real, imag} */,
  {32'h4318d48a, 32'h4194ddea} /* (19, 6, 7) {real, imag} */,
  {32'h3fc7c980, 32'hc115bf18} /* (19, 6, 6) {real, imag} */,
  {32'h42deb268, 32'h419e10b0} /* (19, 6, 5) {real, imag} */,
  {32'hc2281bc0, 32'h3dedc200} /* (19, 6, 4) {real, imag} */,
  {32'hc2922014, 32'h42819ca5} /* (19, 6, 3) {real, imag} */,
  {32'h44538b6f, 32'h4438faac} /* (19, 6, 2) {real, imag} */,
  {32'hc56123f8, 32'hc507f18b} /* (19, 6, 1) {real, imag} */,
  {32'hc57385e8, 32'h00000000} /* (19, 6, 0) {real, imag} */,
  {32'hc558e9f0, 32'h4532516d} /* (19, 5, 31) {real, imag} */,
  {32'h42dab478, 32'hc463ad54} /* (19, 5, 30) {real, imag} */,
  {32'h4289faec, 32'hc31eb606} /* (19, 5, 29) {real, imag} */,
  {32'h4068ef80, 32'hc182aa8c} /* (19, 5, 28) {real, imag} */,
  {32'h43608bab, 32'h42fb30b0} /* (19, 5, 27) {real, imag} */,
  {32'h434813fa, 32'hc2a92f11} /* (19, 5, 26) {real, imag} */,
  {32'hc279c292, 32'h41cb7857} /* (19, 5, 25) {real, imag} */,
  {32'h403a35b0, 32'hc2b4059c} /* (19, 5, 24) {real, imag} */,
  {32'h424189b4, 32'hc1d6f408} /* (19, 5, 23) {real, imag} */,
  {32'h430f3ede, 32'hc1be86ac} /* (19, 5, 22) {real, imag} */,
  {32'h428a48a6, 32'hc2a67ec4} /* (19, 5, 21) {real, imag} */,
  {32'h40edb98e, 32'h4249d398} /* (19, 5, 20) {real, imag} */,
  {32'hc1dd82bc, 32'h41b4f33a} /* (19, 5, 19) {real, imag} */,
  {32'hc18870f3, 32'h42bf1833} /* (19, 5, 18) {real, imag} */,
  {32'hc05495e4, 32'hc2ef6744} /* (19, 5, 17) {real, imag} */,
  {32'h4257eca9, 32'h00000000} /* (19, 5, 16) {real, imag} */,
  {32'hc05495e4, 32'h42ef6744} /* (19, 5, 15) {real, imag} */,
  {32'hc18870f3, 32'hc2bf1833} /* (19, 5, 14) {real, imag} */,
  {32'hc1dd82bc, 32'hc1b4f33a} /* (19, 5, 13) {real, imag} */,
  {32'h40edb98e, 32'hc249d398} /* (19, 5, 12) {real, imag} */,
  {32'h428a48a6, 32'h42a67ec4} /* (19, 5, 11) {real, imag} */,
  {32'h430f3ede, 32'h41be86ac} /* (19, 5, 10) {real, imag} */,
  {32'h424189b4, 32'h41d6f408} /* (19, 5, 9) {real, imag} */,
  {32'h403a35b0, 32'h42b4059c} /* (19, 5, 8) {real, imag} */,
  {32'hc279c292, 32'hc1cb7857} /* (19, 5, 7) {real, imag} */,
  {32'h434813fa, 32'h42a92f11} /* (19, 5, 6) {real, imag} */,
  {32'h43608bab, 32'hc2fb30b0} /* (19, 5, 5) {real, imag} */,
  {32'h4068ef80, 32'h4182aa8c} /* (19, 5, 4) {real, imag} */,
  {32'h4289faec, 32'h431eb606} /* (19, 5, 3) {real, imag} */,
  {32'h42dab478, 32'h4463ad54} /* (19, 5, 2) {real, imag} */,
  {32'hc558e9f0, 32'hc532516d} /* (19, 5, 1) {real, imag} */,
  {32'hc5813d3e, 32'h00000000} /* (19, 5, 0) {real, imag} */,
  {32'hc543fc7c, 32'h455a2266} /* (19, 4, 31) {real, imag} */,
  {32'hc39b0a8e, 32'hc48dce0f} /* (19, 4, 30) {real, imag} */,
  {32'h42c21060, 32'hc233aeb8} /* (19, 4, 29) {real, imag} */,
  {32'h43385d54, 32'hc2a32689} /* (19, 4, 28) {real, imag} */,
  {32'h4373b035, 32'h4342363d} /* (19, 4, 27) {real, imag} */,
  {32'h41c6d9b0, 32'hc1fc7962} /* (19, 4, 26) {real, imag} */,
  {32'h4003c980, 32'h42877eac} /* (19, 4, 25) {real, imag} */,
  {32'hc26d48f6, 32'hc1ec0cb6} /* (19, 4, 24) {real, imag} */,
  {32'h4249ba20, 32'h41c1b78e} /* (19, 4, 23) {real, imag} */,
  {32'h428334d1, 32'hc2573a0f} /* (19, 4, 22) {real, imag} */,
  {32'h42944c40, 32'hc2e0f475} /* (19, 4, 21) {real, imag} */,
  {32'h3f781420, 32'h43122fd4} /* (19, 4, 20) {real, imag} */,
  {32'h4212d1af, 32'h4191e5e1} /* (19, 4, 19) {real, imag} */,
  {32'hc1dfe3c4, 32'hc1d3b144} /* (19, 4, 18) {real, imag} */,
  {32'h423cdb2a, 32'h40d19194} /* (19, 4, 17) {real, imag} */,
  {32'h42fedb80, 32'h00000000} /* (19, 4, 16) {real, imag} */,
  {32'h423cdb2a, 32'hc0d19194} /* (19, 4, 15) {real, imag} */,
  {32'hc1dfe3c4, 32'h41d3b144} /* (19, 4, 14) {real, imag} */,
  {32'h4212d1af, 32'hc191e5e1} /* (19, 4, 13) {real, imag} */,
  {32'h3f781420, 32'hc3122fd4} /* (19, 4, 12) {real, imag} */,
  {32'h42944c40, 32'h42e0f475} /* (19, 4, 11) {real, imag} */,
  {32'h428334d1, 32'h42573a0f} /* (19, 4, 10) {real, imag} */,
  {32'h4249ba20, 32'hc1c1b78e} /* (19, 4, 9) {real, imag} */,
  {32'hc26d48f6, 32'h41ec0cb6} /* (19, 4, 8) {real, imag} */,
  {32'h4003c980, 32'hc2877eac} /* (19, 4, 7) {real, imag} */,
  {32'h41c6d9b0, 32'h41fc7962} /* (19, 4, 6) {real, imag} */,
  {32'h4373b035, 32'hc342363d} /* (19, 4, 5) {real, imag} */,
  {32'h43385d54, 32'h42a32689} /* (19, 4, 4) {real, imag} */,
  {32'h42c21060, 32'h4233aeb8} /* (19, 4, 3) {real, imag} */,
  {32'hc39b0a8e, 32'h448dce0f} /* (19, 4, 2) {real, imag} */,
  {32'hc543fc7c, 32'hc55a2266} /* (19, 4, 1) {real, imag} */,
  {32'hc58d3c0a, 32'h00000000} /* (19, 4, 0) {real, imag} */,
  {32'hc5379e9f, 32'h456ad55a} /* (19, 3, 31) {real, imag} */,
  {32'hc3c5989a, 32'hc4a11b56} /* (19, 3, 30) {real, imag} */,
  {32'h41dc5e69, 32'hc34a646e} /* (19, 3, 29) {real, imag} */,
  {32'h433c6192, 32'hc32d91f0} /* (19, 3, 28) {real, imag} */,
  {32'h43525656, 32'h43280ae3} /* (19, 3, 27) {real, imag} */,
  {32'hc1cdf6b8, 32'h418cfec4} /* (19, 3, 26) {real, imag} */,
  {32'hc288b280, 32'hc295069a} /* (19, 3, 25) {real, imag} */,
  {32'h41b42c9f, 32'hbe679000} /* (19, 3, 24) {real, imag} */,
  {32'h42b96370, 32'hc2ace434} /* (19, 3, 23) {real, imag} */,
  {32'hc239189e, 32'hc249ec9c} /* (19, 3, 22) {real, imag} */,
  {32'h418ac41a, 32'h422856c0} /* (19, 3, 21) {real, imag} */,
  {32'h4147ac54, 32'hc1ec5895} /* (19, 3, 20) {real, imag} */,
  {32'hc157a18b, 32'h42a4e87c} /* (19, 3, 19) {real, imag} */,
  {32'h428963e2, 32'hc182dbdc} /* (19, 3, 18) {real, imag} */,
  {32'hc1b086de, 32'hc02f6d22} /* (19, 3, 17) {real, imag} */,
  {32'hbfaffe80, 32'h00000000} /* (19, 3, 16) {real, imag} */,
  {32'hc1b086de, 32'h402f6d22} /* (19, 3, 15) {real, imag} */,
  {32'h428963e2, 32'h4182dbdc} /* (19, 3, 14) {real, imag} */,
  {32'hc157a18b, 32'hc2a4e87c} /* (19, 3, 13) {real, imag} */,
  {32'h4147ac54, 32'h41ec5895} /* (19, 3, 12) {real, imag} */,
  {32'h418ac41a, 32'hc22856c0} /* (19, 3, 11) {real, imag} */,
  {32'hc239189e, 32'h4249ec9c} /* (19, 3, 10) {real, imag} */,
  {32'h42b96370, 32'h42ace434} /* (19, 3, 9) {real, imag} */,
  {32'h41b42c9f, 32'h3e679000} /* (19, 3, 8) {real, imag} */,
  {32'hc288b280, 32'h4295069a} /* (19, 3, 7) {real, imag} */,
  {32'hc1cdf6b8, 32'hc18cfec4} /* (19, 3, 6) {real, imag} */,
  {32'h43525656, 32'hc3280ae3} /* (19, 3, 5) {real, imag} */,
  {32'h433c6192, 32'h432d91f0} /* (19, 3, 4) {real, imag} */,
  {32'h41dc5e69, 32'h434a646e} /* (19, 3, 3) {real, imag} */,
  {32'hc3c5989a, 32'h44a11b56} /* (19, 3, 2) {real, imag} */,
  {32'hc5379e9f, 32'hc56ad55a} /* (19, 3, 1) {real, imag} */,
  {32'hc58fbc9b, 32'h00000000} /* (19, 3, 0) {real, imag} */,
  {32'hc536a121, 32'h455df71c} /* (19, 2, 31) {real, imag} */,
  {32'hc3e9084c, 32'hc4957f2a} /* (19, 2, 30) {real, imag} */,
  {32'h41f2f560, 32'hc33e8044} /* (19, 2, 29) {real, imag} */,
  {32'h42908872, 32'hc3911941} /* (19, 2, 28) {real, imag} */,
  {32'h436f5eb8, 32'h4367f0f8} /* (19, 2, 27) {real, imag} */,
  {32'h42fb0e83, 32'hc2e24b3b} /* (19, 2, 26) {real, imag} */,
  {32'hc26be798, 32'hc11356fc} /* (19, 2, 25) {real, imag} */,
  {32'h433ba7ae, 32'h430f7ae6} /* (19, 2, 24) {real, imag} */,
  {32'h42abc51c, 32'hc2a74150} /* (19, 2, 23) {real, imag} */,
  {32'h421bcecb, 32'hc2412ce8} /* (19, 2, 22) {real, imag} */,
  {32'h423efff6, 32'h4208325b} /* (19, 2, 21) {real, imag} */,
  {32'h42380c9b, 32'hc232d332} /* (19, 2, 20) {real, imag} */,
  {32'hc290dd38, 32'hc2de107c} /* (19, 2, 19) {real, imag} */,
  {32'h41313114, 32'h416fe0aa} /* (19, 2, 18) {real, imag} */,
  {32'h40d187a4, 32'h41c53a3a} /* (19, 2, 17) {real, imag} */,
  {32'hc10f347c, 32'h00000000} /* (19, 2, 16) {real, imag} */,
  {32'h40d187a4, 32'hc1c53a3a} /* (19, 2, 15) {real, imag} */,
  {32'h41313114, 32'hc16fe0aa} /* (19, 2, 14) {real, imag} */,
  {32'hc290dd38, 32'h42de107c} /* (19, 2, 13) {real, imag} */,
  {32'h42380c9b, 32'h4232d332} /* (19, 2, 12) {real, imag} */,
  {32'h423efff6, 32'hc208325b} /* (19, 2, 11) {real, imag} */,
  {32'h421bcecb, 32'h42412ce8} /* (19, 2, 10) {real, imag} */,
  {32'h42abc51c, 32'h42a74150} /* (19, 2, 9) {real, imag} */,
  {32'h433ba7ae, 32'hc30f7ae6} /* (19, 2, 8) {real, imag} */,
  {32'hc26be798, 32'h411356fc} /* (19, 2, 7) {real, imag} */,
  {32'h42fb0e83, 32'h42e24b3b} /* (19, 2, 6) {real, imag} */,
  {32'h436f5eb8, 32'hc367f0f8} /* (19, 2, 5) {real, imag} */,
  {32'h42908872, 32'h43911941} /* (19, 2, 4) {real, imag} */,
  {32'h41f2f560, 32'h433e8044} /* (19, 2, 3) {real, imag} */,
  {32'hc3e9084c, 32'h44957f2a} /* (19, 2, 2) {real, imag} */,
  {32'hc536a121, 32'hc55df71c} /* (19, 2, 1) {real, imag} */,
  {32'hc596af9f, 32'h00000000} /* (19, 2, 0) {real, imag} */,
  {32'hc5422d01, 32'h454b56be} /* (19, 1, 31) {real, imag} */,
  {32'hc3946f6d, 32'hc47c0826} /* (19, 1, 30) {real, imag} */,
  {32'h42d82def, 32'hc2b211c8} /* (19, 1, 29) {real, imag} */,
  {32'h42af613e, 32'hc3953ef6} /* (19, 1, 28) {real, imag} */,
  {32'h4354e030, 32'h42cd7aff} /* (19, 1, 27) {real, imag} */,
  {32'h430b5df5, 32'hc34a3f4c} /* (19, 1, 26) {real, imag} */,
  {32'hc20482be, 32'h43151b5a} /* (19, 1, 25) {real, imag} */,
  {32'h4173ccf8, 32'hc24a10c6} /* (19, 1, 24) {real, imag} */,
  {32'hc2345bd6, 32'h4263cd96} /* (19, 1, 23) {real, imag} */,
  {32'hc28a81f5, 32'hc267deea} /* (19, 1, 22) {real, imag} */,
  {32'hc2af594e, 32'h40989fe4} /* (19, 1, 21) {real, imag} */,
  {32'h4202541a, 32'hc2424c50} /* (19, 1, 20) {real, imag} */,
  {32'h4233da3c, 32'hc21b4c0a} /* (19, 1, 19) {real, imag} */,
  {32'h4243f24a, 32'hc1df8965} /* (19, 1, 18) {real, imag} */,
  {32'h40ffb6a9, 32'h41f27f23} /* (19, 1, 17) {real, imag} */,
  {32'h420bc4c1, 32'h00000000} /* (19, 1, 16) {real, imag} */,
  {32'h40ffb6a9, 32'hc1f27f23} /* (19, 1, 15) {real, imag} */,
  {32'h4243f24a, 32'h41df8965} /* (19, 1, 14) {real, imag} */,
  {32'h4233da3c, 32'h421b4c0a} /* (19, 1, 13) {real, imag} */,
  {32'h4202541a, 32'h42424c50} /* (19, 1, 12) {real, imag} */,
  {32'hc2af594e, 32'hc0989fe4} /* (19, 1, 11) {real, imag} */,
  {32'hc28a81f5, 32'h4267deea} /* (19, 1, 10) {real, imag} */,
  {32'hc2345bd6, 32'hc263cd96} /* (19, 1, 9) {real, imag} */,
  {32'h4173ccf8, 32'h424a10c6} /* (19, 1, 8) {real, imag} */,
  {32'hc20482be, 32'hc3151b5a} /* (19, 1, 7) {real, imag} */,
  {32'h430b5df5, 32'h434a3f4c} /* (19, 1, 6) {real, imag} */,
  {32'h4354e030, 32'hc2cd7aff} /* (19, 1, 5) {real, imag} */,
  {32'h42af613e, 32'h43953ef6} /* (19, 1, 4) {real, imag} */,
  {32'h42d82def, 32'h42b211c8} /* (19, 1, 3) {real, imag} */,
  {32'hc3946f6d, 32'h447c0826} /* (19, 1, 2) {real, imag} */,
  {32'hc5422d01, 32'hc54b56be} /* (19, 1, 1) {real, imag} */,
  {32'hc597a309, 32'h00000000} /* (19, 1, 0) {real, imag} */,
  {32'hc55214c8, 32'h4527e45c} /* (19, 0, 31) {real, imag} */,
  {32'h42b064c0, 32'hc43ad0f4} /* (19, 0, 30) {real, imag} */,
  {32'h425c66e9, 32'hc260dc5e} /* (19, 0, 29) {real, imag} */,
  {32'h41d19244, 32'hc2ea71e8} /* (19, 0, 28) {real, imag} */,
  {32'h4239446c, 32'h421397a6} /* (19, 0, 27) {real, imag} */,
  {32'h41e5a90e, 32'h4151b11a} /* (19, 0, 26) {real, imag} */,
  {32'hc1eebe82, 32'h4263b6de} /* (19, 0, 25) {real, imag} */,
  {32'hc2a81c08, 32'hc25080b0} /* (19, 0, 24) {real, imag} */,
  {32'hc2074f35, 32'h410f6d04} /* (19, 0, 23) {real, imag} */,
  {32'h410d469c, 32'h40a7adc0} /* (19, 0, 22) {real, imag} */,
  {32'h42132eae, 32'h41d6ffcc} /* (19, 0, 21) {real, imag} */,
  {32'h40e852e4, 32'hc1073574} /* (19, 0, 20) {real, imag} */,
  {32'h418d3a22, 32'h401a98e0} /* (19, 0, 19) {real, imag} */,
  {32'h421722aa, 32'hc29b7a99} /* (19, 0, 18) {real, imag} */,
  {32'h4232dd56, 32'hc1b26d43} /* (19, 0, 17) {real, imag} */,
  {32'h4260bc9a, 32'h00000000} /* (19, 0, 16) {real, imag} */,
  {32'h4232dd56, 32'h41b26d43} /* (19, 0, 15) {real, imag} */,
  {32'h421722aa, 32'h429b7a99} /* (19, 0, 14) {real, imag} */,
  {32'h418d3a22, 32'hc01a98e0} /* (19, 0, 13) {real, imag} */,
  {32'h40e852e4, 32'h41073574} /* (19, 0, 12) {real, imag} */,
  {32'h42132eae, 32'hc1d6ffcc} /* (19, 0, 11) {real, imag} */,
  {32'h410d469c, 32'hc0a7adc0} /* (19, 0, 10) {real, imag} */,
  {32'hc2074f35, 32'hc10f6d04} /* (19, 0, 9) {real, imag} */,
  {32'hc2a81c08, 32'h425080b0} /* (19, 0, 8) {real, imag} */,
  {32'hc1eebe82, 32'hc263b6de} /* (19, 0, 7) {real, imag} */,
  {32'h41e5a90e, 32'hc151b11a} /* (19, 0, 6) {real, imag} */,
  {32'h4239446c, 32'hc21397a6} /* (19, 0, 5) {real, imag} */,
  {32'h41d19244, 32'h42ea71e8} /* (19, 0, 4) {real, imag} */,
  {32'h425c66e9, 32'h4260dc5e} /* (19, 0, 3) {real, imag} */,
  {32'h42b064c0, 32'h443ad0f4} /* (19, 0, 2) {real, imag} */,
  {32'hc55214c8, 32'hc527e45c} /* (19, 0, 1) {real, imag} */,
  {32'hc5907501, 32'h00000000} /* (19, 0, 0) {real, imag} */,
  {32'hc5485909, 32'h44cd20fe} /* (18, 31, 31) {real, imag} */,
  {32'h441271f9, 32'hc3f38109} /* (18, 31, 30) {real, imag} */,
  {32'h42ba7b6b, 32'h42a948ba} /* (18, 31, 29) {real, imag} */,
  {32'hc1c7dad9, 32'hc22250da} /* (18, 31, 28) {real, imag} */,
  {32'h427a7fa2, 32'hc2b5a1ca} /* (18, 31, 27) {real, imag} */,
  {32'h42b42166, 32'h3ff498f0} /* (18, 31, 26) {real, imag} */,
  {32'h4223d509, 32'h423a506e} /* (18, 31, 25) {real, imag} */,
  {32'hc2195e25, 32'hc22f5376} /* (18, 31, 24) {real, imag} */,
  {32'h42583b66, 32'hc2465e42} /* (18, 31, 23) {real, imag} */,
  {32'hc1d7f8a1, 32'h4292aaeb} /* (18, 31, 22) {real, imag} */,
  {32'hc19927f6, 32'h42aaaf50} /* (18, 31, 21) {real, imag} */,
  {32'hc291b142, 32'hc0dfde88} /* (18, 31, 20) {real, imag} */,
  {32'hc23cd29a, 32'hc2783bbe} /* (18, 31, 19) {real, imag} */,
  {32'hc0e04298, 32'hc29245a2} /* (18, 31, 18) {real, imag} */,
  {32'h420dbbb2, 32'h41583d56} /* (18, 31, 17) {real, imag} */,
  {32'h421e888c, 32'h00000000} /* (18, 31, 16) {real, imag} */,
  {32'h420dbbb2, 32'hc1583d56} /* (18, 31, 15) {real, imag} */,
  {32'hc0e04298, 32'h429245a2} /* (18, 31, 14) {real, imag} */,
  {32'hc23cd29a, 32'h42783bbe} /* (18, 31, 13) {real, imag} */,
  {32'hc291b142, 32'h40dfde88} /* (18, 31, 12) {real, imag} */,
  {32'hc19927f6, 32'hc2aaaf50} /* (18, 31, 11) {real, imag} */,
  {32'hc1d7f8a1, 32'hc292aaeb} /* (18, 31, 10) {real, imag} */,
  {32'h42583b66, 32'h42465e42} /* (18, 31, 9) {real, imag} */,
  {32'hc2195e25, 32'h422f5376} /* (18, 31, 8) {real, imag} */,
  {32'h4223d509, 32'hc23a506e} /* (18, 31, 7) {real, imag} */,
  {32'h42b42166, 32'hbff498f0} /* (18, 31, 6) {real, imag} */,
  {32'h427a7fa2, 32'h42b5a1ca} /* (18, 31, 5) {real, imag} */,
  {32'hc1c7dad9, 32'h422250da} /* (18, 31, 4) {real, imag} */,
  {32'h42ba7b6b, 32'hc2a948ba} /* (18, 31, 3) {real, imag} */,
  {32'h441271f9, 32'h43f38109} /* (18, 31, 2) {real, imag} */,
  {32'hc5485909, 32'hc4cd20fe} /* (18, 31, 1) {real, imag} */,
  {32'hc575da3e, 32'h00000000} /* (18, 31, 0) {real, imag} */,
  {32'hc57420a4, 32'h44b46214} /* (18, 30, 31) {real, imag} */,
  {32'h4475fd44, 32'hc3c8ebf0} /* (18, 30, 30) {real, imag} */,
  {32'h42c69b41, 32'h435a41e3} /* (18, 30, 29) {real, imag} */,
  {32'hc2c97f33, 32'h4206de40} /* (18, 30, 28) {real, imag} */,
  {32'h4351f0e8, 32'hc2ca790b} /* (18, 30, 27) {real, imag} */,
  {32'h422da416, 32'h40cfd876} /* (18, 30, 26) {real, imag} */,
  {32'h425ff5b2, 32'h430f1f64} /* (18, 30, 25) {real, imag} */,
  {32'h426782a8, 32'hc2ad3ff6} /* (18, 30, 24) {real, imag} */,
  {32'h423f9596, 32'hc285e9d2} /* (18, 30, 23) {real, imag} */,
  {32'hc1be06a0, 32'h42908893} /* (18, 30, 22) {real, imag} */,
  {32'hc271b85d, 32'hc29ff154} /* (18, 30, 21) {real, imag} */,
  {32'hc2555374, 32'h411294d4} /* (18, 30, 20) {real, imag} */,
  {32'h42fcd8be, 32'h42c03eb2} /* (18, 30, 19) {real, imag} */,
  {32'h42bf950a, 32'h429d9e82} /* (18, 30, 18) {real, imag} */,
  {32'h41b9196e, 32'h419e6a75} /* (18, 30, 17) {real, imag} */,
  {32'hc26d8676, 32'h00000000} /* (18, 30, 16) {real, imag} */,
  {32'h41b9196e, 32'hc19e6a75} /* (18, 30, 15) {real, imag} */,
  {32'h42bf950a, 32'hc29d9e82} /* (18, 30, 14) {real, imag} */,
  {32'h42fcd8be, 32'hc2c03eb2} /* (18, 30, 13) {real, imag} */,
  {32'hc2555374, 32'hc11294d4} /* (18, 30, 12) {real, imag} */,
  {32'hc271b85d, 32'h429ff154} /* (18, 30, 11) {real, imag} */,
  {32'hc1be06a0, 32'hc2908893} /* (18, 30, 10) {real, imag} */,
  {32'h423f9596, 32'h4285e9d2} /* (18, 30, 9) {real, imag} */,
  {32'h426782a8, 32'h42ad3ff6} /* (18, 30, 8) {real, imag} */,
  {32'h425ff5b2, 32'hc30f1f64} /* (18, 30, 7) {real, imag} */,
  {32'h422da416, 32'hc0cfd876} /* (18, 30, 6) {real, imag} */,
  {32'h4351f0e8, 32'h42ca790b} /* (18, 30, 5) {real, imag} */,
  {32'hc2c97f33, 32'hc206de40} /* (18, 30, 4) {real, imag} */,
  {32'h42c69b41, 32'hc35a41e3} /* (18, 30, 3) {real, imag} */,
  {32'h4475fd44, 32'h43c8ebf0} /* (18, 30, 2) {real, imag} */,
  {32'hc57420a4, 32'hc4b46214} /* (18, 30, 1) {real, imag} */,
  {32'hc57b8391, 32'h00000000} /* (18, 30, 0) {real, imag} */,
  {32'hc581b6ac, 32'h448af024} /* (18, 29, 31) {real, imag} */,
  {32'h4498a024, 32'hc3dceb3e} /* (18, 29, 30) {real, imag} */,
  {32'h3fc3b2c0, 32'h423c1039} /* (18, 29, 29) {real, imag} */,
  {32'hc3231138, 32'h42f45228} /* (18, 29, 28) {real, imag} */,
  {32'h42c52f29, 32'h41e40ab4} /* (18, 29, 27) {real, imag} */,
  {32'h43279f4c, 32'h42934cd2} /* (18, 29, 26) {real, imag} */,
  {32'h41973c95, 32'h42de25da} /* (18, 29, 25) {real, imag} */,
  {32'h41df70df, 32'h4116e826} /* (18, 29, 24) {real, imag} */,
  {32'hc3075cc7, 32'hc20a7bd5} /* (18, 29, 23) {real, imag} */,
  {32'h41e1bf26, 32'hc2a8ae9b} /* (18, 29, 22) {real, imag} */,
  {32'hc2527046, 32'hc2c56f68} /* (18, 29, 21) {real, imag} */,
  {32'hc27ec09d, 32'hc24fac4a} /* (18, 29, 20) {real, imag} */,
  {32'hc1162eea, 32'hc192b87f} /* (18, 29, 19) {real, imag} */,
  {32'h3f3d66c8, 32'hc28754ee} /* (18, 29, 18) {real, imag} */,
  {32'hc0d80fbc, 32'h41b263a6} /* (18, 29, 17) {real, imag} */,
  {32'h41b6b657, 32'h00000000} /* (18, 29, 16) {real, imag} */,
  {32'hc0d80fbc, 32'hc1b263a6} /* (18, 29, 15) {real, imag} */,
  {32'h3f3d66c8, 32'h428754ee} /* (18, 29, 14) {real, imag} */,
  {32'hc1162eea, 32'h4192b87f} /* (18, 29, 13) {real, imag} */,
  {32'hc27ec09d, 32'h424fac4a} /* (18, 29, 12) {real, imag} */,
  {32'hc2527046, 32'h42c56f68} /* (18, 29, 11) {real, imag} */,
  {32'h41e1bf26, 32'h42a8ae9b} /* (18, 29, 10) {real, imag} */,
  {32'hc3075cc7, 32'h420a7bd5} /* (18, 29, 9) {real, imag} */,
  {32'h41df70df, 32'hc116e826} /* (18, 29, 8) {real, imag} */,
  {32'h41973c95, 32'hc2de25da} /* (18, 29, 7) {real, imag} */,
  {32'h43279f4c, 32'hc2934cd2} /* (18, 29, 6) {real, imag} */,
  {32'h42c52f29, 32'hc1e40ab4} /* (18, 29, 5) {real, imag} */,
  {32'hc3231138, 32'hc2f45228} /* (18, 29, 4) {real, imag} */,
  {32'h3fc3b2c0, 32'hc23c1039} /* (18, 29, 3) {real, imag} */,
  {32'h4498a024, 32'h43dceb3e} /* (18, 29, 2) {real, imag} */,
  {32'hc581b6ac, 32'hc48af024} /* (18, 29, 1) {real, imag} */,
  {32'hc57e2241, 32'h00000000} /* (18, 29, 0) {real, imag} */,
  {32'hc584f7a1, 32'h44764337} /* (18, 28, 31) {real, imag} */,
  {32'h44b80218, 32'hc3fb5fc4} /* (18, 28, 30) {real, imag} */,
  {32'h40fda580, 32'hc2697808} /* (18, 28, 29) {real, imag} */,
  {32'hc36c614b, 32'h42d260d8} /* (18, 28, 28) {real, imag} */,
  {32'h428b8d82, 32'hc249c079} /* (18, 28, 27) {real, imag} */,
  {32'h42fc5082, 32'h40b95f74} /* (18, 28, 26) {real, imag} */,
  {32'hc2104c32, 32'hc2f2398a} /* (18, 28, 25) {real, imag} */,
  {32'hc0f46cdc, 32'hc2d1a35f} /* (18, 28, 24) {real, imag} */,
  {32'hc198246c, 32'h42f28c1c} /* (18, 28, 23) {real, imag} */,
  {32'hc2b5f1ca, 32'h41cea5ea} /* (18, 28, 22) {real, imag} */,
  {32'h42608428, 32'hc29c11ee} /* (18, 28, 21) {real, imag} */,
  {32'hc05cfc94, 32'h412bef64} /* (18, 28, 20) {real, imag} */,
  {32'hc248261e, 32'h4021f7d0} /* (18, 28, 19) {real, imag} */,
  {32'hc1074b9c, 32'hc2064eb2} /* (18, 28, 18) {real, imag} */,
  {32'hc1d030ff, 32'hc09b24b0} /* (18, 28, 17) {real, imag} */,
  {32'h4104fbcc, 32'h00000000} /* (18, 28, 16) {real, imag} */,
  {32'hc1d030ff, 32'h409b24b0} /* (18, 28, 15) {real, imag} */,
  {32'hc1074b9c, 32'h42064eb2} /* (18, 28, 14) {real, imag} */,
  {32'hc248261e, 32'hc021f7d0} /* (18, 28, 13) {real, imag} */,
  {32'hc05cfc94, 32'hc12bef64} /* (18, 28, 12) {real, imag} */,
  {32'h42608428, 32'h429c11ee} /* (18, 28, 11) {real, imag} */,
  {32'hc2b5f1ca, 32'hc1cea5ea} /* (18, 28, 10) {real, imag} */,
  {32'hc198246c, 32'hc2f28c1c} /* (18, 28, 9) {real, imag} */,
  {32'hc0f46cdc, 32'h42d1a35f} /* (18, 28, 8) {real, imag} */,
  {32'hc2104c32, 32'h42f2398a} /* (18, 28, 7) {real, imag} */,
  {32'h42fc5082, 32'hc0b95f74} /* (18, 28, 6) {real, imag} */,
  {32'h428b8d82, 32'h4249c079} /* (18, 28, 5) {real, imag} */,
  {32'hc36c614b, 32'hc2d260d8} /* (18, 28, 4) {real, imag} */,
  {32'h40fda580, 32'h42697808} /* (18, 28, 3) {real, imag} */,
  {32'h44b80218, 32'h43fb5fc4} /* (18, 28, 2) {real, imag} */,
  {32'hc584f7a1, 32'hc4764337} /* (18, 28, 1) {real, imag} */,
  {32'hc581e0fa, 32'h00000000} /* (18, 28, 0) {real, imag} */,
  {32'hc58429df, 32'h4428df60} /* (18, 27, 31) {real, imag} */,
  {32'h44bf1e69, 32'hc4048e8a} /* (18, 27, 30) {real, imag} */,
  {32'h421b2b12, 32'hc1b72595} /* (18, 27, 29) {real, imag} */,
  {32'hc35a7d90, 32'hc21a921e} /* (18, 27, 28) {real, imag} */,
  {32'h42b7cd00, 32'h41643ad4} /* (18, 27, 27) {real, imag} */,
  {32'hc25da1e0, 32'h42d4785e} /* (18, 27, 26) {real, imag} */,
  {32'h408d7cac, 32'hc1865142} /* (18, 27, 25) {real, imag} */,
  {32'hc1976db7, 32'hc2db4484} /* (18, 27, 24) {real, imag} */,
  {32'h41abea79, 32'hc2c947ce} /* (18, 27, 23) {real, imag} */,
  {32'hc1e8078a, 32'h41876187} /* (18, 27, 22) {real, imag} */,
  {32'h426b72eb, 32'hc29933d4} /* (18, 27, 21) {real, imag} */,
  {32'h42b4beaa, 32'h4240036c} /* (18, 27, 20) {real, imag} */,
  {32'h416d3b8a, 32'hc21e8303} /* (18, 27, 19) {real, imag} */,
  {32'h422c46a4, 32'hc2058394} /* (18, 27, 18) {real, imag} */,
  {32'hc10ec83e, 32'hc19c8f2d} /* (18, 27, 17) {real, imag} */,
  {32'h41a6f2dc, 32'h00000000} /* (18, 27, 16) {real, imag} */,
  {32'hc10ec83e, 32'h419c8f2d} /* (18, 27, 15) {real, imag} */,
  {32'h422c46a4, 32'h42058394} /* (18, 27, 14) {real, imag} */,
  {32'h416d3b8a, 32'h421e8303} /* (18, 27, 13) {real, imag} */,
  {32'h42b4beaa, 32'hc240036c} /* (18, 27, 12) {real, imag} */,
  {32'h426b72eb, 32'h429933d4} /* (18, 27, 11) {real, imag} */,
  {32'hc1e8078a, 32'hc1876187} /* (18, 27, 10) {real, imag} */,
  {32'h41abea79, 32'h42c947ce} /* (18, 27, 9) {real, imag} */,
  {32'hc1976db7, 32'h42db4484} /* (18, 27, 8) {real, imag} */,
  {32'h408d7cac, 32'h41865142} /* (18, 27, 7) {real, imag} */,
  {32'hc25da1e0, 32'hc2d4785e} /* (18, 27, 6) {real, imag} */,
  {32'h42b7cd00, 32'hc1643ad4} /* (18, 27, 5) {real, imag} */,
  {32'hc35a7d90, 32'h421a921e} /* (18, 27, 4) {real, imag} */,
  {32'h421b2b12, 32'h41b72595} /* (18, 27, 3) {real, imag} */,
  {32'h44bf1e69, 32'h44048e8a} /* (18, 27, 2) {real, imag} */,
  {32'hc58429df, 32'hc428df60} /* (18, 27, 1) {real, imag} */,
  {32'hc581594d, 32'h00000000} /* (18, 27, 0) {real, imag} */,
  {32'hc57dcd48, 32'h4407282c} /* (18, 26, 31) {real, imag} */,
  {32'h44b2d5e9, 32'hc40f3042} /* (18, 26, 30) {real, imag} */,
  {32'hc2233766, 32'hc20e6d82} /* (18, 26, 29) {real, imag} */,
  {32'hc3898ac8, 32'hc2893597} /* (18, 26, 28) {real, imag} */,
  {32'h42ce28f2, 32'hc1fa29ae} /* (18, 26, 27) {real, imag} */,
  {32'h41b70e2d, 32'h4281fe06} /* (18, 26, 26) {real, imag} */,
  {32'h41d42cec, 32'h409a6dc4} /* (18, 26, 25) {real, imag} */,
  {32'h42451530, 32'hc2e32530} /* (18, 26, 24) {real, imag} */,
  {32'hc1f93996, 32'hc28ad9f6} /* (18, 26, 23) {real, imag} */,
  {32'h429fa1de, 32'hc1bfcc56} /* (18, 26, 22) {real, imag} */,
  {32'h424226e2, 32'h418a424d} /* (18, 26, 21) {real, imag} */,
  {32'h427744a3, 32'h42366ed0} /* (18, 26, 20) {real, imag} */,
  {32'hc2b54612, 32'hc236315e} /* (18, 26, 19) {real, imag} */,
  {32'h42b08157, 32'hc2332cb6} /* (18, 26, 18) {real, imag} */,
  {32'hc21e07a1, 32'h3f76d6c0} /* (18, 26, 17) {real, imag} */,
  {32'h421d1152, 32'h00000000} /* (18, 26, 16) {real, imag} */,
  {32'hc21e07a1, 32'hbf76d6c0} /* (18, 26, 15) {real, imag} */,
  {32'h42b08157, 32'h42332cb6} /* (18, 26, 14) {real, imag} */,
  {32'hc2b54612, 32'h4236315e} /* (18, 26, 13) {real, imag} */,
  {32'h427744a3, 32'hc2366ed0} /* (18, 26, 12) {real, imag} */,
  {32'h424226e2, 32'hc18a424d} /* (18, 26, 11) {real, imag} */,
  {32'h429fa1de, 32'h41bfcc56} /* (18, 26, 10) {real, imag} */,
  {32'hc1f93996, 32'h428ad9f6} /* (18, 26, 9) {real, imag} */,
  {32'h42451530, 32'h42e32530} /* (18, 26, 8) {real, imag} */,
  {32'h41d42cec, 32'hc09a6dc4} /* (18, 26, 7) {real, imag} */,
  {32'h41b70e2d, 32'hc281fe06} /* (18, 26, 6) {real, imag} */,
  {32'h42ce28f2, 32'h41fa29ae} /* (18, 26, 5) {real, imag} */,
  {32'hc3898ac8, 32'h42893597} /* (18, 26, 4) {real, imag} */,
  {32'hc2233766, 32'h420e6d82} /* (18, 26, 3) {real, imag} */,
  {32'h44b2d5e9, 32'h440f3042} /* (18, 26, 2) {real, imag} */,
  {32'hc57dcd48, 32'hc407282c} /* (18, 26, 1) {real, imag} */,
  {32'hc5806fe4, 32'h00000000} /* (18, 26, 0) {real, imag} */,
  {32'hc56d031c, 32'h43d63550} /* (18, 25, 31) {real, imag} */,
  {32'h44ae8b52, 32'hc3815ce8} /* (18, 25, 30) {real, imag} */,
  {32'h429e27c2, 32'hc26d72f1} /* (18, 25, 29) {real, imag} */,
  {32'hc3d19550, 32'hc2aa2bb8} /* (18, 25, 28) {real, imag} */,
  {32'h43718903, 32'hc3858523} /* (18, 25, 27) {real, imag} */,
  {32'hc2e5ae0c, 32'hc2681d47} /* (18, 25, 26) {real, imag} */,
  {32'hc1e537d8, 32'h4348df32} /* (18, 25, 25) {real, imag} */,
  {32'h4315cc26, 32'hc2e33ff1} /* (18, 25, 24) {real, imag} */,
  {32'hc29b6b1f, 32'h4268c9f6} /* (18, 25, 23) {real, imag} */,
  {32'h4300da9b, 32'hc3117666} /* (18, 25, 22) {real, imag} */,
  {32'hc21b14c1, 32'hc2d765b3} /* (18, 25, 21) {real, imag} */,
  {32'hc25a0de9, 32'h43394612} /* (18, 25, 20) {real, imag} */,
  {32'h42b36809, 32'hc2a15c27} /* (18, 25, 19) {real, imag} */,
  {32'h416f905c, 32'h4186dd74} /* (18, 25, 18) {real, imag} */,
  {32'h4122831a, 32'h41abdcb4} /* (18, 25, 17) {real, imag} */,
  {32'h42c41d80, 32'h00000000} /* (18, 25, 16) {real, imag} */,
  {32'h4122831a, 32'hc1abdcb4} /* (18, 25, 15) {real, imag} */,
  {32'h416f905c, 32'hc186dd74} /* (18, 25, 14) {real, imag} */,
  {32'h42b36809, 32'h42a15c27} /* (18, 25, 13) {real, imag} */,
  {32'hc25a0de9, 32'hc3394612} /* (18, 25, 12) {real, imag} */,
  {32'hc21b14c1, 32'h42d765b3} /* (18, 25, 11) {real, imag} */,
  {32'h4300da9b, 32'h43117666} /* (18, 25, 10) {real, imag} */,
  {32'hc29b6b1f, 32'hc268c9f6} /* (18, 25, 9) {real, imag} */,
  {32'h4315cc26, 32'h42e33ff1} /* (18, 25, 8) {real, imag} */,
  {32'hc1e537d8, 32'hc348df32} /* (18, 25, 7) {real, imag} */,
  {32'hc2e5ae0c, 32'h42681d47} /* (18, 25, 6) {real, imag} */,
  {32'h43718903, 32'h43858523} /* (18, 25, 5) {real, imag} */,
  {32'hc3d19550, 32'h42aa2bb8} /* (18, 25, 4) {real, imag} */,
  {32'h429e27c2, 32'h426d72f1} /* (18, 25, 3) {real, imag} */,
  {32'h44ae8b52, 32'h43815ce8} /* (18, 25, 2) {real, imag} */,
  {32'hc56d031c, 32'hc3d63550} /* (18, 25, 1) {real, imag} */,
  {32'hc56b02bc, 32'h00000000} /* (18, 25, 0) {real, imag} */,
  {32'hc54e023e, 32'h4381a1c8} /* (18, 24, 31) {real, imag} */,
  {32'h44a2c872, 32'hc31b0720} /* (18, 24, 30) {real, imag} */,
  {32'hc04fc8d0, 32'hc2eb1202} /* (18, 24, 29) {real, imag} */,
  {32'hc3a4f64b, 32'hc1d247f4} /* (18, 24, 28) {real, imag} */,
  {32'h43859b66, 32'hc3284f00} /* (18, 24, 27) {real, imag} */,
  {32'hc28ab50c, 32'hc2b9ecc8} /* (18, 24, 26) {real, imag} */,
  {32'hc0fc6798, 32'h42d71060} /* (18, 24, 25) {real, imag} */,
  {32'h42ba11eb, 32'hc21ca4aa} /* (18, 24, 24) {real, imag} */,
  {32'hc2c30f30, 32'hbf6d0770} /* (18, 24, 23) {real, imag} */,
  {32'h417e0d90, 32'h420a6ad2} /* (18, 24, 22) {real, imag} */,
  {32'h41b456a8, 32'hc2dc36fe} /* (18, 24, 21) {real, imag} */,
  {32'h429c4b04, 32'h4281a9c4} /* (18, 24, 20) {real, imag} */,
  {32'h424c7434, 32'h422d5766} /* (18, 24, 19) {real, imag} */,
  {32'h41eac914, 32'hc237ab1b} /* (18, 24, 18) {real, imag} */,
  {32'h425983bc, 32'hc161e479} /* (18, 24, 17) {real, imag} */,
  {32'hc2a8d139, 32'h00000000} /* (18, 24, 16) {real, imag} */,
  {32'h425983bc, 32'h4161e479} /* (18, 24, 15) {real, imag} */,
  {32'h41eac914, 32'h4237ab1b} /* (18, 24, 14) {real, imag} */,
  {32'h424c7434, 32'hc22d5766} /* (18, 24, 13) {real, imag} */,
  {32'h429c4b04, 32'hc281a9c4} /* (18, 24, 12) {real, imag} */,
  {32'h41b456a8, 32'h42dc36fe} /* (18, 24, 11) {real, imag} */,
  {32'h417e0d90, 32'hc20a6ad2} /* (18, 24, 10) {real, imag} */,
  {32'hc2c30f30, 32'h3f6d0770} /* (18, 24, 9) {real, imag} */,
  {32'h42ba11eb, 32'h421ca4aa} /* (18, 24, 8) {real, imag} */,
  {32'hc0fc6798, 32'hc2d71060} /* (18, 24, 7) {real, imag} */,
  {32'hc28ab50c, 32'h42b9ecc8} /* (18, 24, 6) {real, imag} */,
  {32'h43859b66, 32'h43284f00} /* (18, 24, 5) {real, imag} */,
  {32'hc3a4f64b, 32'h41d247f4} /* (18, 24, 4) {real, imag} */,
  {32'hc04fc8d0, 32'h42eb1202} /* (18, 24, 3) {real, imag} */,
  {32'h44a2c872, 32'h431b0720} /* (18, 24, 2) {real, imag} */,
  {32'hc54e023e, 32'hc381a1c8} /* (18, 24, 1) {real, imag} */,
  {32'hc55568d0, 32'h00000000} /* (18, 24, 0) {real, imag} */,
  {32'hc52c152a, 32'h43547600} /* (18, 23, 31) {real, imag} */,
  {32'h4491b6d8, 32'hc33c5cdc} /* (18, 23, 30) {real, imag} */,
  {32'hc2e52a56, 32'hc3007e8b} /* (18, 23, 29) {real, imag} */,
  {32'hc323a7d6, 32'hc24b4228} /* (18, 23, 28) {real, imag} */,
  {32'h4381d14a, 32'hc3112f15} /* (18, 23, 27) {real, imag} */,
  {32'h42b45d4e, 32'hc2850af5} /* (18, 23, 26) {real, imag} */,
  {32'hc29fd136, 32'hc2160803} /* (18, 23, 25) {real, imag} */,
  {32'h42e8a390, 32'h40e8fe50} /* (18, 23, 24) {real, imag} */,
  {32'hc2da3ec1, 32'h420b4763} /* (18, 23, 23) {real, imag} */,
  {32'h41bc459e, 32'h4269c690} /* (18, 23, 22) {real, imag} */,
  {32'h42bf4250, 32'hc25caf4c} /* (18, 23, 21) {real, imag} */,
  {32'hc1c4dfb6, 32'h42057f5a} /* (18, 23, 20) {real, imag} */,
  {32'h4191c4bc, 32'h42077514} /* (18, 23, 19) {real, imag} */,
  {32'h40a4bd8c, 32'h410cb596} /* (18, 23, 18) {real, imag} */,
  {32'hc1c9700e, 32'hc1f30e84} /* (18, 23, 17) {real, imag} */,
  {32'hc29f2a8d, 32'h00000000} /* (18, 23, 16) {real, imag} */,
  {32'hc1c9700e, 32'h41f30e84} /* (18, 23, 15) {real, imag} */,
  {32'h40a4bd8c, 32'hc10cb596} /* (18, 23, 14) {real, imag} */,
  {32'h4191c4bc, 32'hc2077514} /* (18, 23, 13) {real, imag} */,
  {32'hc1c4dfb6, 32'hc2057f5a} /* (18, 23, 12) {real, imag} */,
  {32'h42bf4250, 32'h425caf4c} /* (18, 23, 11) {real, imag} */,
  {32'h41bc459e, 32'hc269c690} /* (18, 23, 10) {real, imag} */,
  {32'hc2da3ec1, 32'hc20b4763} /* (18, 23, 9) {real, imag} */,
  {32'h42e8a390, 32'hc0e8fe50} /* (18, 23, 8) {real, imag} */,
  {32'hc29fd136, 32'h42160803} /* (18, 23, 7) {real, imag} */,
  {32'h42b45d4e, 32'h42850af5} /* (18, 23, 6) {real, imag} */,
  {32'h4381d14a, 32'h43112f15} /* (18, 23, 5) {real, imag} */,
  {32'hc323a7d6, 32'h424b4228} /* (18, 23, 4) {real, imag} */,
  {32'hc2e52a56, 32'h43007e8b} /* (18, 23, 3) {real, imag} */,
  {32'h4491b6d8, 32'h433c5cdc} /* (18, 23, 2) {real, imag} */,
  {32'hc52c152a, 32'hc3547600} /* (18, 23, 1) {real, imag} */,
  {32'hc52d7d72, 32'h00000000} /* (18, 23, 0) {real, imag} */,
  {32'hc4f92926, 32'h432caabe} /* (18, 22, 31) {real, imag} */,
  {32'h446643bd, 32'hc1fe2d80} /* (18, 22, 30) {real, imag} */,
  {32'hc3295874, 32'h421064bd} /* (18, 22, 29) {real, imag} */,
  {32'hc1396dc8, 32'h42239474} /* (18, 22, 28) {real, imag} */,
  {32'h42f4131d, 32'hc343e0b4} /* (18, 22, 27) {real, imag} */,
  {32'hc20811aa, 32'hc2f6d140} /* (18, 22, 26) {real, imag} */,
  {32'hc31d7913, 32'hc2436959} /* (18, 22, 25) {real, imag} */,
  {32'h409c6c64, 32'h42ae8a30} /* (18, 22, 24) {real, imag} */,
  {32'h4129f4c0, 32'hbfcbca20} /* (18, 22, 23) {real, imag} */,
  {32'h418a00cf, 32'hc237ca14} /* (18, 22, 22) {real, imag} */,
  {32'h41a15da9, 32'h412292b8} /* (18, 22, 21) {real, imag} */,
  {32'hc207d70b, 32'h4218f3f6} /* (18, 22, 20) {real, imag} */,
  {32'h42007c55, 32'hc29700ce} /* (18, 22, 19) {real, imag} */,
  {32'h41a0683b, 32'hc10a7d4a} /* (18, 22, 18) {real, imag} */,
  {32'hc12653c8, 32'hc24e98d1} /* (18, 22, 17) {real, imag} */,
  {32'h42163652, 32'h00000000} /* (18, 22, 16) {real, imag} */,
  {32'hc12653c8, 32'h424e98d1} /* (18, 22, 15) {real, imag} */,
  {32'h41a0683b, 32'h410a7d4a} /* (18, 22, 14) {real, imag} */,
  {32'h42007c55, 32'h429700ce} /* (18, 22, 13) {real, imag} */,
  {32'hc207d70b, 32'hc218f3f6} /* (18, 22, 12) {real, imag} */,
  {32'h41a15da9, 32'hc12292b8} /* (18, 22, 11) {real, imag} */,
  {32'h418a00cf, 32'h4237ca14} /* (18, 22, 10) {real, imag} */,
  {32'h4129f4c0, 32'h3fcbca20} /* (18, 22, 9) {real, imag} */,
  {32'h409c6c64, 32'hc2ae8a30} /* (18, 22, 8) {real, imag} */,
  {32'hc31d7913, 32'h42436959} /* (18, 22, 7) {real, imag} */,
  {32'hc20811aa, 32'h42f6d140} /* (18, 22, 6) {real, imag} */,
  {32'h42f4131d, 32'h4343e0b4} /* (18, 22, 5) {real, imag} */,
  {32'hc1396dc8, 32'hc2239474} /* (18, 22, 4) {real, imag} */,
  {32'hc3295874, 32'hc21064bd} /* (18, 22, 3) {real, imag} */,
  {32'h446643bd, 32'h41fe2d80} /* (18, 22, 2) {real, imag} */,
  {32'hc4f92926, 32'hc32caabe} /* (18, 22, 1) {real, imag} */,
  {32'hc5034fe4, 32'h00000000} /* (18, 22, 0) {real, imag} */,
  {32'hc440a4bb, 32'h4318d112} /* (18, 21, 31) {real, imag} */,
  {32'h4399ce8e, 32'h430634ae} /* (18, 21, 30) {real, imag} */,
  {32'hc2b1785a, 32'h421b0220} /* (18, 21, 29) {real, imag} */,
  {32'hc1bca76a, 32'h423b7c7a} /* (18, 21, 28) {real, imag} */,
  {32'h4274c374, 32'hc2ebe66e} /* (18, 21, 27) {real, imag} */,
  {32'hc25cfe1a, 32'h41bb0956} /* (18, 21, 26) {real, imag} */,
  {32'h4254aea2, 32'h4292c276} /* (18, 21, 25) {real, imag} */,
  {32'h42883785, 32'hc25f77ac} /* (18, 21, 24) {real, imag} */,
  {32'h422076f8, 32'hc2101fcc} /* (18, 21, 23) {real, imag} */,
  {32'h42a9e936, 32'hc29945f7} /* (18, 21, 22) {real, imag} */,
  {32'h41a42be0, 32'hc2aa2bfb} /* (18, 21, 21) {real, imag} */,
  {32'h424d2e90, 32'h3e7c4280} /* (18, 21, 20) {real, imag} */,
  {32'h411e75a2, 32'h41610305} /* (18, 21, 19) {real, imag} */,
  {32'hc1cbbecc, 32'hc134f4b0} /* (18, 21, 18) {real, imag} */,
  {32'h40577d58, 32'h41939ba8} /* (18, 21, 17) {real, imag} */,
  {32'h40cd8ca6, 32'h00000000} /* (18, 21, 16) {real, imag} */,
  {32'h40577d58, 32'hc1939ba8} /* (18, 21, 15) {real, imag} */,
  {32'hc1cbbecc, 32'h4134f4b0} /* (18, 21, 14) {real, imag} */,
  {32'h411e75a2, 32'hc1610305} /* (18, 21, 13) {real, imag} */,
  {32'h424d2e90, 32'hbe7c4280} /* (18, 21, 12) {real, imag} */,
  {32'h41a42be0, 32'h42aa2bfb} /* (18, 21, 11) {real, imag} */,
  {32'h42a9e936, 32'h429945f7} /* (18, 21, 10) {real, imag} */,
  {32'h422076f8, 32'h42101fcc} /* (18, 21, 9) {real, imag} */,
  {32'h42883785, 32'h425f77ac} /* (18, 21, 8) {real, imag} */,
  {32'h4254aea2, 32'hc292c276} /* (18, 21, 7) {real, imag} */,
  {32'hc25cfe1a, 32'hc1bb0956} /* (18, 21, 6) {real, imag} */,
  {32'h4274c374, 32'h42ebe66e} /* (18, 21, 5) {real, imag} */,
  {32'hc1bca76a, 32'hc23b7c7a} /* (18, 21, 4) {real, imag} */,
  {32'hc2b1785a, 32'hc21b0220} /* (18, 21, 3) {real, imag} */,
  {32'h4399ce8e, 32'hc30634ae} /* (18, 21, 2) {real, imag} */,
  {32'hc440a4bb, 32'hc318d112} /* (18, 21, 1) {real, imag} */,
  {32'hc494b6f6, 32'h00000000} /* (18, 21, 0) {real, imag} */,
  {32'h445d2809, 32'hc198e660} /* (18, 20, 31) {real, imag} */,
  {32'hc3bf33f6, 32'h43a2ba84} /* (18, 20, 30) {real, imag} */,
  {32'hc1644590, 32'h41a95ab4} /* (18, 20, 29) {real, imag} */,
  {32'h436670fd, 32'h41c4629b} /* (18, 20, 28) {real, imag} */,
  {32'hc2c4ef9c, 32'h42b2d91b} /* (18, 20, 27) {real, imag} */,
  {32'hc30ec652, 32'h4276cccf} /* (18, 20, 26) {real, imag} */,
  {32'h430f5fa0, 32'hc29218ce} /* (18, 20, 25) {real, imag} */,
  {32'h42052613, 32'hc2bf5ed8} /* (18, 20, 24) {real, imag} */,
  {32'hc17a02d8, 32'h4163fa6a} /* (18, 20, 23) {real, imag} */,
  {32'h420bb436, 32'h41d2800d} /* (18, 20, 22) {real, imag} */,
  {32'hc257dbd4, 32'hc1ae3fa8} /* (18, 20, 21) {real, imag} */,
  {32'hc21f98de, 32'hc23c76c4} /* (18, 20, 20) {real, imag} */,
  {32'h42b9564c, 32'h406b0f60} /* (18, 20, 19) {real, imag} */,
  {32'hc18676a6, 32'h42398fa9} /* (18, 20, 18) {real, imag} */,
  {32'h425a2cb2, 32'hc232c01d} /* (18, 20, 17) {real, imag} */,
  {32'hc14b7870, 32'h00000000} /* (18, 20, 16) {real, imag} */,
  {32'h425a2cb2, 32'h4232c01d} /* (18, 20, 15) {real, imag} */,
  {32'hc18676a6, 32'hc2398fa9} /* (18, 20, 14) {real, imag} */,
  {32'h42b9564c, 32'hc06b0f60} /* (18, 20, 13) {real, imag} */,
  {32'hc21f98de, 32'h423c76c4} /* (18, 20, 12) {real, imag} */,
  {32'hc257dbd4, 32'h41ae3fa8} /* (18, 20, 11) {real, imag} */,
  {32'h420bb436, 32'hc1d2800d} /* (18, 20, 10) {real, imag} */,
  {32'hc17a02d8, 32'hc163fa6a} /* (18, 20, 9) {real, imag} */,
  {32'h42052613, 32'h42bf5ed8} /* (18, 20, 8) {real, imag} */,
  {32'h430f5fa0, 32'h429218ce} /* (18, 20, 7) {real, imag} */,
  {32'hc30ec652, 32'hc276cccf} /* (18, 20, 6) {real, imag} */,
  {32'hc2c4ef9c, 32'hc2b2d91b} /* (18, 20, 5) {real, imag} */,
  {32'h436670fd, 32'hc1c4629b} /* (18, 20, 4) {real, imag} */,
  {32'hc1644590, 32'hc1a95ab4} /* (18, 20, 3) {real, imag} */,
  {32'hc3bf33f6, 32'hc3a2ba84} /* (18, 20, 2) {real, imag} */,
  {32'h445d2809, 32'h4198e660} /* (18, 20, 1) {real, imag} */,
  {32'h431848bc, 32'h00000000} /* (18, 20, 0) {real, imag} */,
  {32'h44fc919e, 32'hc2f6050c} /* (18, 19, 31) {real, imag} */,
  {32'hc44dfd48, 32'h438b66fa} /* (18, 19, 30) {real, imag} */,
  {32'hc1d09e60, 32'h42802130} /* (18, 19, 29) {real, imag} */,
  {32'h43bb2050, 32'hc2877edf} /* (18, 19, 28) {real, imag} */,
  {32'hc300d0ec, 32'h43068c87} /* (18, 19, 27) {real, imag} */,
  {32'hc33a8ea1, 32'h42cd0b53} /* (18, 19, 26) {real, imag} */,
  {32'h423c0cb7, 32'hc1e7ae12} /* (18, 19, 25) {real, imag} */,
  {32'hc0ee6214, 32'h425e2d44} /* (18, 19, 24) {real, imag} */,
  {32'hc12dc722, 32'h428058e3} /* (18, 19, 23) {real, imag} */,
  {32'hc28dd71e, 32'hc29d759c} /* (18, 19, 22) {real, imag} */,
  {32'hc2e8a810, 32'h42e9cae3} /* (18, 19, 21) {real, imag} */,
  {32'h416a88db, 32'hc201513a} /* (18, 19, 20) {real, imag} */,
  {32'hc28d975e, 32'hc2aeae05} /* (18, 19, 19) {real, imag} */,
  {32'h4112a635, 32'h41ea7988} /* (18, 19, 18) {real, imag} */,
  {32'hc0091800, 32'h41ae8af6} /* (18, 19, 17) {real, imag} */,
  {32'h425312ea, 32'h00000000} /* (18, 19, 16) {real, imag} */,
  {32'hc0091800, 32'hc1ae8af6} /* (18, 19, 15) {real, imag} */,
  {32'h4112a635, 32'hc1ea7988} /* (18, 19, 14) {real, imag} */,
  {32'hc28d975e, 32'h42aeae05} /* (18, 19, 13) {real, imag} */,
  {32'h416a88db, 32'h4201513a} /* (18, 19, 12) {real, imag} */,
  {32'hc2e8a810, 32'hc2e9cae3} /* (18, 19, 11) {real, imag} */,
  {32'hc28dd71e, 32'h429d759c} /* (18, 19, 10) {real, imag} */,
  {32'hc12dc722, 32'hc28058e3} /* (18, 19, 9) {real, imag} */,
  {32'hc0ee6214, 32'hc25e2d44} /* (18, 19, 8) {real, imag} */,
  {32'h423c0cb7, 32'h41e7ae12} /* (18, 19, 7) {real, imag} */,
  {32'hc33a8ea1, 32'hc2cd0b53} /* (18, 19, 6) {real, imag} */,
  {32'hc300d0ec, 32'hc3068c87} /* (18, 19, 5) {real, imag} */,
  {32'h43bb2050, 32'h42877edf} /* (18, 19, 4) {real, imag} */,
  {32'hc1d09e60, 32'hc2802130} /* (18, 19, 3) {real, imag} */,
  {32'hc44dfd48, 32'hc38b66fa} /* (18, 19, 2) {real, imag} */,
  {32'h44fc919e, 32'h42f6050c} /* (18, 19, 1) {real, imag} */,
  {32'h449a844a, 32'h00000000} /* (18, 19, 0) {real, imag} */,
  {32'h452e6a4d, 32'hc38f5a98} /* (18, 18, 31) {real, imag} */,
  {32'hc487dfd6, 32'h432dd2f3} /* (18, 18, 30) {real, imag} */,
  {32'h42b50537, 32'hc2cf8424} /* (18, 18, 29) {real, imag} */,
  {32'h43ca0803, 32'hc30509be} /* (18, 18, 28) {real, imag} */,
  {32'hc31b5b90, 32'h42dbfb1a} /* (18, 18, 27) {real, imag} */,
  {32'hc2f47c71, 32'hc216e156} /* (18, 18, 26) {real, imag} */,
  {32'h419a3ea2, 32'hc1f342dc} /* (18, 18, 25) {real, imag} */,
  {32'hc0b2959c, 32'h4204c33a} /* (18, 18, 24) {real, imag} */,
  {32'hc1836308, 32'h428a8e98} /* (18, 18, 23) {real, imag} */,
  {32'hc27b2d4d, 32'h41f7aa85} /* (18, 18, 22) {real, imag} */,
  {32'hc2791703, 32'h422c0e68} /* (18, 18, 21) {real, imag} */,
  {32'hc1e5d630, 32'h42b56018} /* (18, 18, 20) {real, imag} */,
  {32'hc22cb096, 32'h41d60f65} /* (18, 18, 19) {real, imag} */,
  {32'h415c5cf6, 32'h417dcf95} /* (18, 18, 18) {real, imag} */,
  {32'hc02a7ce0, 32'h41f4edd8} /* (18, 18, 17) {real, imag} */,
  {32'hc227c0ff, 32'h00000000} /* (18, 18, 16) {real, imag} */,
  {32'hc02a7ce0, 32'hc1f4edd8} /* (18, 18, 15) {real, imag} */,
  {32'h415c5cf6, 32'hc17dcf95} /* (18, 18, 14) {real, imag} */,
  {32'hc22cb096, 32'hc1d60f65} /* (18, 18, 13) {real, imag} */,
  {32'hc1e5d630, 32'hc2b56018} /* (18, 18, 12) {real, imag} */,
  {32'hc2791703, 32'hc22c0e68} /* (18, 18, 11) {real, imag} */,
  {32'hc27b2d4d, 32'hc1f7aa85} /* (18, 18, 10) {real, imag} */,
  {32'hc1836308, 32'hc28a8e98} /* (18, 18, 9) {real, imag} */,
  {32'hc0b2959c, 32'hc204c33a} /* (18, 18, 8) {real, imag} */,
  {32'h419a3ea2, 32'h41f342dc} /* (18, 18, 7) {real, imag} */,
  {32'hc2f47c71, 32'h4216e156} /* (18, 18, 6) {real, imag} */,
  {32'hc31b5b90, 32'hc2dbfb1a} /* (18, 18, 5) {real, imag} */,
  {32'h43ca0803, 32'h430509be} /* (18, 18, 4) {real, imag} */,
  {32'h42b50537, 32'h42cf8424} /* (18, 18, 3) {real, imag} */,
  {32'hc487dfd6, 32'hc32dd2f3} /* (18, 18, 2) {real, imag} */,
  {32'h452e6a4d, 32'h438f5a98} /* (18, 18, 1) {real, imag} */,
  {32'h44e3b4de, 32'h00000000} /* (18, 18, 0) {real, imag} */,
  {32'h4548b463, 32'hc38bc34d} /* (18, 17, 31) {real, imag} */,
  {32'hc498d860, 32'h432f7f82} /* (18, 17, 30) {real, imag} */,
  {32'h42ae050f, 32'hc2dda6ae} /* (18, 17, 29) {real, imag} */,
  {32'h43aafa66, 32'hc23a063a} /* (18, 17, 28) {real, imag} */,
  {32'hc3853773, 32'h43021b1c} /* (18, 17, 27) {real, imag} */,
  {32'hc25b0054, 32'hc135642c} /* (18, 17, 26) {real, imag} */,
  {32'h430e2973, 32'hc1c0862f} /* (18, 17, 25) {real, imag} */,
  {32'hc2cd9d11, 32'h40d3b11e} /* (18, 17, 24) {real, imag} */,
  {32'hc1d42e23, 32'hc2bd635a} /* (18, 17, 23) {real, imag} */,
  {32'h4220905b, 32'hc1c821a0} /* (18, 17, 22) {real, imag} */,
  {32'hbfe5a188, 32'h4237202e} /* (18, 17, 21) {real, imag} */,
  {32'h41e1054f, 32'hc1337489} /* (18, 17, 20) {real, imag} */,
  {32'hc20e639e, 32'h4295bad9} /* (18, 17, 19) {real, imag} */,
  {32'h42a1547d, 32'hc2134890} /* (18, 17, 18) {real, imag} */,
  {32'h4268300d, 32'hc1df0b3c} /* (18, 17, 17) {real, imag} */,
  {32'hc0b56fe3, 32'h00000000} /* (18, 17, 16) {real, imag} */,
  {32'h4268300d, 32'h41df0b3c} /* (18, 17, 15) {real, imag} */,
  {32'h42a1547d, 32'h42134890} /* (18, 17, 14) {real, imag} */,
  {32'hc20e639e, 32'hc295bad9} /* (18, 17, 13) {real, imag} */,
  {32'h41e1054f, 32'h41337489} /* (18, 17, 12) {real, imag} */,
  {32'hbfe5a188, 32'hc237202e} /* (18, 17, 11) {real, imag} */,
  {32'h4220905b, 32'h41c821a0} /* (18, 17, 10) {real, imag} */,
  {32'hc1d42e23, 32'h42bd635a} /* (18, 17, 9) {real, imag} */,
  {32'hc2cd9d11, 32'hc0d3b11e} /* (18, 17, 8) {real, imag} */,
  {32'h430e2973, 32'h41c0862f} /* (18, 17, 7) {real, imag} */,
  {32'hc25b0054, 32'h4135642c} /* (18, 17, 6) {real, imag} */,
  {32'hc3853773, 32'hc3021b1c} /* (18, 17, 5) {real, imag} */,
  {32'h43aafa66, 32'h423a063a} /* (18, 17, 4) {real, imag} */,
  {32'h42ae050f, 32'h42dda6ae} /* (18, 17, 3) {real, imag} */,
  {32'hc498d860, 32'hc32f7f82} /* (18, 17, 2) {real, imag} */,
  {32'h4548b463, 32'h438bc34d} /* (18, 17, 1) {real, imag} */,
  {32'h45089bae, 32'h00000000} /* (18, 17, 0) {real, imag} */,
  {32'h455761b8, 32'hc38511e0} /* (18, 16, 31) {real, imag} */,
  {32'hc4bcb132, 32'h426aac00} /* (18, 16, 30) {real, imag} */,
  {32'h42c402fe, 32'hc2984ce6} /* (18, 16, 29) {real, imag} */,
  {32'h43a1f033, 32'h4203b72e} /* (18, 16, 28) {real, imag} */,
  {32'hc3a58dd0, 32'h430d5af1} /* (18, 16, 27) {real, imag} */,
  {32'hc27ac634, 32'h4240802f} /* (18, 16, 26) {real, imag} */,
  {32'h426adc82, 32'hc232a59a} /* (18, 16, 25) {real, imag} */,
  {32'hc2db7e2e, 32'h42cd7c1c} /* (18, 16, 24) {real, imag} */,
  {32'hc1825a6e, 32'h423aa93e} /* (18, 16, 23) {real, imag} */,
  {32'hc29aadd2, 32'h42ae2cdb} /* (18, 16, 22) {real, imag} */,
  {32'hbecf9e20, 32'h428d3f80} /* (18, 16, 21) {real, imag} */,
  {32'h431a4785, 32'hc1dfe39f} /* (18, 16, 20) {real, imag} */,
  {32'hc27dae2a, 32'h3f3c1c70} /* (18, 16, 19) {real, imag} */,
  {32'hc2267a0f, 32'h41c07c14} /* (18, 16, 18) {real, imag} */,
  {32'h41968668, 32'hc1c94128} /* (18, 16, 17) {real, imag} */,
  {32'hc2f19f17, 32'h00000000} /* (18, 16, 16) {real, imag} */,
  {32'h41968668, 32'h41c94128} /* (18, 16, 15) {real, imag} */,
  {32'hc2267a0f, 32'hc1c07c14} /* (18, 16, 14) {real, imag} */,
  {32'hc27dae2a, 32'hbf3c1c70} /* (18, 16, 13) {real, imag} */,
  {32'h431a4785, 32'h41dfe39f} /* (18, 16, 12) {real, imag} */,
  {32'hbecf9e20, 32'hc28d3f80} /* (18, 16, 11) {real, imag} */,
  {32'hc29aadd2, 32'hc2ae2cdb} /* (18, 16, 10) {real, imag} */,
  {32'hc1825a6e, 32'hc23aa93e} /* (18, 16, 9) {real, imag} */,
  {32'hc2db7e2e, 32'hc2cd7c1c} /* (18, 16, 8) {real, imag} */,
  {32'h426adc82, 32'h4232a59a} /* (18, 16, 7) {real, imag} */,
  {32'hc27ac634, 32'hc240802f} /* (18, 16, 6) {real, imag} */,
  {32'hc3a58dd0, 32'hc30d5af1} /* (18, 16, 5) {real, imag} */,
  {32'h43a1f033, 32'hc203b72e} /* (18, 16, 4) {real, imag} */,
  {32'h42c402fe, 32'h42984ce6} /* (18, 16, 3) {real, imag} */,
  {32'hc4bcb132, 32'hc26aac00} /* (18, 16, 2) {real, imag} */,
  {32'h455761b8, 32'h438511e0} /* (18, 16, 1) {real, imag} */,
  {32'h451d93aa, 32'h00000000} /* (18, 16, 0) {real, imag} */,
  {32'h45566965, 32'hc39feacb} /* (18, 15, 31) {real, imag} */,
  {32'hc4be4800, 32'h439c3d48} /* (18, 15, 30) {real, imag} */,
  {32'h42e8710d, 32'hc2d4929e} /* (18, 15, 29) {real, imag} */,
  {32'h435294cb, 32'hc17bdf18} /* (18, 15, 28) {real, imag} */,
  {32'hc32d9c58, 32'h438727c7} /* (18, 15, 27) {real, imag} */,
  {32'h41707340, 32'hc0f7e130} /* (18, 15, 26) {real, imag} */,
  {32'h41163130, 32'hc238cd66} /* (18, 15, 25) {real, imag} */,
  {32'h422b99c2, 32'h4219038c} /* (18, 15, 24) {real, imag} */,
  {32'h42abe40d, 32'h4209668c} /* (18, 15, 23) {real, imag} */,
  {32'h4263f605, 32'h430d970c} /* (18, 15, 22) {real, imag} */,
  {32'hc17531bf, 32'h43361964} /* (18, 15, 21) {real, imag} */,
  {32'h41cbf2cf, 32'h406b6f74} /* (18, 15, 20) {real, imag} */,
  {32'h41a27e83, 32'hc188ad5f} /* (18, 15, 19) {real, imag} */,
  {32'hc251063e, 32'h420c8c62} /* (18, 15, 18) {real, imag} */,
  {32'hc1ea7fc6, 32'h426ddf2a} /* (18, 15, 17) {real, imag} */,
  {32'h410b6784, 32'h00000000} /* (18, 15, 16) {real, imag} */,
  {32'hc1ea7fc6, 32'hc26ddf2a} /* (18, 15, 15) {real, imag} */,
  {32'hc251063e, 32'hc20c8c62} /* (18, 15, 14) {real, imag} */,
  {32'h41a27e83, 32'h4188ad5f} /* (18, 15, 13) {real, imag} */,
  {32'h41cbf2cf, 32'hc06b6f74} /* (18, 15, 12) {real, imag} */,
  {32'hc17531bf, 32'hc3361964} /* (18, 15, 11) {real, imag} */,
  {32'h4263f605, 32'hc30d970c} /* (18, 15, 10) {real, imag} */,
  {32'h42abe40d, 32'hc209668c} /* (18, 15, 9) {real, imag} */,
  {32'h422b99c2, 32'hc219038c} /* (18, 15, 8) {real, imag} */,
  {32'h41163130, 32'h4238cd66} /* (18, 15, 7) {real, imag} */,
  {32'h41707340, 32'h40f7e130} /* (18, 15, 6) {real, imag} */,
  {32'hc32d9c58, 32'hc38727c7} /* (18, 15, 5) {real, imag} */,
  {32'h435294cb, 32'h417bdf18} /* (18, 15, 4) {real, imag} */,
  {32'h42e8710d, 32'h42d4929e} /* (18, 15, 3) {real, imag} */,
  {32'hc4be4800, 32'hc39c3d48} /* (18, 15, 2) {real, imag} */,
  {32'h45566965, 32'h439feacb} /* (18, 15, 1) {real, imag} */,
  {32'h4519da1a, 32'h00000000} /* (18, 15, 0) {real, imag} */,
  {32'h4540d2a7, 32'hc3387150} /* (18, 14, 31) {real, imag} */,
  {32'hc4af9f82, 32'h43acfa1e} /* (18, 14, 30) {real, imag} */,
  {32'h437d7a1a, 32'hc2f7a7fc} /* (18, 14, 29) {real, imag} */,
  {32'h4355f65a, 32'hc0c27130} /* (18, 14, 28) {real, imag} */,
  {32'hc37b85e8, 32'h4377059b} /* (18, 14, 27) {real, imag} */,
  {32'h42fc1d5f, 32'h425748c2} /* (18, 14, 26) {real, imag} */,
  {32'hc299a45e, 32'hc299dc36} /* (18, 14, 25) {real, imag} */,
  {32'hc1f88eed, 32'h42df7633} /* (18, 14, 24) {real, imag} */,
  {32'hc2554c60, 32'h42929298} /* (18, 14, 23) {real, imag} */,
  {32'h428379b1, 32'hc2aa8153} /* (18, 14, 22) {real, imag} */,
  {32'hc201040f, 32'h42146ed4} /* (18, 14, 21) {real, imag} */,
  {32'hc144ec8d, 32'hc11386a4} /* (18, 14, 20) {real, imag} */,
  {32'hc07cf308, 32'hc28b4bac} /* (18, 14, 19) {real, imag} */,
  {32'hc28519d7, 32'h414287ed} /* (18, 14, 18) {real, imag} */,
  {32'h42166d2c, 32'hbfae01d8} /* (18, 14, 17) {real, imag} */,
  {32'h41aadbda, 32'h00000000} /* (18, 14, 16) {real, imag} */,
  {32'h42166d2c, 32'h3fae01d8} /* (18, 14, 15) {real, imag} */,
  {32'hc28519d7, 32'hc14287ed} /* (18, 14, 14) {real, imag} */,
  {32'hc07cf308, 32'h428b4bac} /* (18, 14, 13) {real, imag} */,
  {32'hc144ec8d, 32'h411386a4} /* (18, 14, 12) {real, imag} */,
  {32'hc201040f, 32'hc2146ed4} /* (18, 14, 11) {real, imag} */,
  {32'h428379b1, 32'h42aa8153} /* (18, 14, 10) {real, imag} */,
  {32'hc2554c60, 32'hc2929298} /* (18, 14, 9) {real, imag} */,
  {32'hc1f88eed, 32'hc2df7633} /* (18, 14, 8) {real, imag} */,
  {32'hc299a45e, 32'h4299dc36} /* (18, 14, 7) {real, imag} */,
  {32'h42fc1d5f, 32'hc25748c2} /* (18, 14, 6) {real, imag} */,
  {32'hc37b85e8, 32'hc377059b} /* (18, 14, 5) {real, imag} */,
  {32'h4355f65a, 32'h40c27130} /* (18, 14, 4) {real, imag} */,
  {32'h437d7a1a, 32'h42f7a7fc} /* (18, 14, 3) {real, imag} */,
  {32'hc4af9f82, 32'hc3acfa1e} /* (18, 14, 2) {real, imag} */,
  {32'h4540d2a7, 32'h43387150} /* (18, 14, 1) {real, imag} */,
  {32'h450f9b89, 32'h00000000} /* (18, 14, 0) {real, imag} */,
  {32'h45256e97, 32'h425ea118} /* (18, 13, 31) {real, imag} */,
  {32'hc4991ee8, 32'h4376802b} /* (18, 13, 30) {real, imag} */,
  {32'h43440f78, 32'hc2a78f4a} /* (18, 13, 29) {real, imag} */,
  {32'h42b5b066, 32'h421a4816} /* (18, 13, 28) {real, imag} */,
  {32'hc3411b8e, 32'h428e1cea} /* (18, 13, 27) {real, imag} */,
  {32'h415928c0, 32'h42de7317} /* (18, 13, 26) {real, imag} */,
  {32'hc229a48b, 32'hc1124d3c} /* (18, 13, 25) {real, imag} */,
  {32'hc287278f, 32'h421224d2} /* (18, 13, 24) {real, imag} */,
  {32'h4263dfc6, 32'h42627fcf} /* (18, 13, 23) {real, imag} */,
  {32'hc1f96de0, 32'hc29215e0} /* (18, 13, 22) {real, imag} */,
  {32'h4063aac0, 32'h424d838a} /* (18, 13, 21) {real, imag} */,
  {32'h420c5783, 32'hc25519fa} /* (18, 13, 20) {real, imag} */,
  {32'h41a95377, 32'h42fe9551} /* (18, 13, 19) {real, imag} */,
  {32'hc1597d1b, 32'h422937a4} /* (18, 13, 18) {real, imag} */,
  {32'h415ac886, 32'h426da5cb} /* (18, 13, 17) {real, imag} */,
  {32'hc2730c2e, 32'h00000000} /* (18, 13, 16) {real, imag} */,
  {32'h415ac886, 32'hc26da5cb} /* (18, 13, 15) {real, imag} */,
  {32'hc1597d1b, 32'hc22937a4} /* (18, 13, 14) {real, imag} */,
  {32'h41a95377, 32'hc2fe9551} /* (18, 13, 13) {real, imag} */,
  {32'h420c5783, 32'h425519fa} /* (18, 13, 12) {real, imag} */,
  {32'h4063aac0, 32'hc24d838a} /* (18, 13, 11) {real, imag} */,
  {32'hc1f96de0, 32'h429215e0} /* (18, 13, 10) {real, imag} */,
  {32'h4263dfc6, 32'hc2627fcf} /* (18, 13, 9) {real, imag} */,
  {32'hc287278f, 32'hc21224d2} /* (18, 13, 8) {real, imag} */,
  {32'hc229a48b, 32'h41124d3c} /* (18, 13, 7) {real, imag} */,
  {32'h415928c0, 32'hc2de7317} /* (18, 13, 6) {real, imag} */,
  {32'hc3411b8e, 32'hc28e1cea} /* (18, 13, 5) {real, imag} */,
  {32'h42b5b066, 32'hc21a4816} /* (18, 13, 4) {real, imag} */,
  {32'h43440f78, 32'h42a78f4a} /* (18, 13, 3) {real, imag} */,
  {32'hc4991ee8, 32'hc376802b} /* (18, 13, 2) {real, imag} */,
  {32'h45256e97, 32'hc25ea118} /* (18, 13, 1) {real, imag} */,
  {32'h44f5599e, 32'h00000000} /* (18, 13, 0) {real, imag} */,
  {32'h44f77e12, 32'h43385a4c} /* (18, 12, 31) {real, imag} */,
  {32'hc47d76f5, 32'h4391d79e} /* (18, 12, 30) {real, imag} */,
  {32'h42c5c33c, 32'hc31a8b8a} /* (18, 12, 29) {real, imag} */,
  {32'h42a1226a, 32'hc2a4750a} /* (18, 12, 28) {real, imag} */,
  {32'hc2e2c7ce, 32'h4305a52a} /* (18, 12, 27) {real, imag} */,
  {32'h42837200, 32'h42266d3b} /* (18, 12, 26) {real, imag} */,
  {32'h42120098, 32'hc2b1256e} /* (18, 12, 25) {real, imag} */,
  {32'hc2103c59, 32'h40e1e4e0} /* (18, 12, 24) {real, imag} */,
  {32'h428b5f4d, 32'hc1f3a34b} /* (18, 12, 23) {real, imag} */,
  {32'h421ef0c0, 32'h41ff966d} /* (18, 12, 22) {real, imag} */,
  {32'h428327f6, 32'h42898033} /* (18, 12, 21) {real, imag} */,
  {32'hc2211bca, 32'hc1cdfedd} /* (18, 12, 20) {real, imag} */,
  {32'h428ea538, 32'h42940567} /* (18, 12, 19) {real, imag} */,
  {32'h42039707, 32'h4259efe7} /* (18, 12, 18) {real, imag} */,
  {32'hc281aa56, 32'h41a7f0de} /* (18, 12, 17) {real, imag} */,
  {32'hc163f928, 32'h00000000} /* (18, 12, 16) {real, imag} */,
  {32'hc281aa56, 32'hc1a7f0de} /* (18, 12, 15) {real, imag} */,
  {32'h42039707, 32'hc259efe7} /* (18, 12, 14) {real, imag} */,
  {32'h428ea538, 32'hc2940567} /* (18, 12, 13) {real, imag} */,
  {32'hc2211bca, 32'h41cdfedd} /* (18, 12, 12) {real, imag} */,
  {32'h428327f6, 32'hc2898033} /* (18, 12, 11) {real, imag} */,
  {32'h421ef0c0, 32'hc1ff966d} /* (18, 12, 10) {real, imag} */,
  {32'h428b5f4d, 32'h41f3a34b} /* (18, 12, 9) {real, imag} */,
  {32'hc2103c59, 32'hc0e1e4e0} /* (18, 12, 8) {real, imag} */,
  {32'h42120098, 32'h42b1256e} /* (18, 12, 7) {real, imag} */,
  {32'h42837200, 32'hc2266d3b} /* (18, 12, 6) {real, imag} */,
  {32'hc2e2c7ce, 32'hc305a52a} /* (18, 12, 5) {real, imag} */,
  {32'h42a1226a, 32'h42a4750a} /* (18, 12, 4) {real, imag} */,
  {32'h42c5c33c, 32'h431a8b8a} /* (18, 12, 3) {real, imag} */,
  {32'hc47d76f5, 32'hc391d79e} /* (18, 12, 2) {real, imag} */,
  {32'h44f77e12, 32'hc3385a4c} /* (18, 12, 1) {real, imag} */,
  {32'h44ac2308, 32'h00000000} /* (18, 12, 0) {real, imag} */,
  {32'h446120db, 32'h43c4f407} /* (18, 11, 31) {real, imag} */,
  {32'hc4135d16, 32'h4347c4e2} /* (18, 11, 30) {real, imag} */,
  {32'h4317cfff, 32'hc1d0965f} /* (18, 11, 29) {real, imag} */,
  {32'h42abfaaa, 32'hc252e246} /* (18, 11, 28) {real, imag} */,
  {32'hc30d0edb, 32'h41b24b18} /* (18, 11, 27) {real, imag} */,
  {32'h42b7ddab, 32'h42fdce14} /* (18, 11, 26) {real, imag} */,
  {32'hc27c9a28, 32'h41dd6262} /* (18, 11, 25) {real, imag} */,
  {32'hc27e98f6, 32'h421a9f24} /* (18, 11, 24) {real, imag} */,
  {32'hc20b0362, 32'h4265a01c} /* (18, 11, 23) {real, imag} */,
  {32'h40c02ee8, 32'hc2c79151} /* (18, 11, 22) {real, imag} */,
  {32'hc2e4eb10, 32'h42df1691} /* (18, 11, 21) {real, imag} */,
  {32'hc2f02620, 32'hc263fde0} /* (18, 11, 20) {real, imag} */,
  {32'h408026b4, 32'h41693451} /* (18, 11, 19) {real, imag} */,
  {32'hc1aae252, 32'h42381d50} /* (18, 11, 18) {real, imag} */,
  {32'h423596ee, 32'hc22e0766} /* (18, 11, 17) {real, imag} */,
  {32'h41dcd068, 32'h00000000} /* (18, 11, 16) {real, imag} */,
  {32'h423596ee, 32'h422e0766} /* (18, 11, 15) {real, imag} */,
  {32'hc1aae252, 32'hc2381d50} /* (18, 11, 14) {real, imag} */,
  {32'h408026b4, 32'hc1693451} /* (18, 11, 13) {real, imag} */,
  {32'hc2f02620, 32'h4263fde0} /* (18, 11, 12) {real, imag} */,
  {32'hc2e4eb10, 32'hc2df1691} /* (18, 11, 11) {real, imag} */,
  {32'h40c02ee8, 32'h42c79151} /* (18, 11, 10) {real, imag} */,
  {32'hc20b0362, 32'hc265a01c} /* (18, 11, 9) {real, imag} */,
  {32'hc27e98f6, 32'hc21a9f24} /* (18, 11, 8) {real, imag} */,
  {32'hc27c9a28, 32'hc1dd6262} /* (18, 11, 7) {real, imag} */,
  {32'h42b7ddab, 32'hc2fdce14} /* (18, 11, 6) {real, imag} */,
  {32'hc30d0edb, 32'hc1b24b18} /* (18, 11, 5) {real, imag} */,
  {32'h42abfaaa, 32'h4252e246} /* (18, 11, 4) {real, imag} */,
  {32'h4317cfff, 32'h41d0965f} /* (18, 11, 3) {real, imag} */,
  {32'hc4135d16, 32'hc347c4e2} /* (18, 11, 2) {real, imag} */,
  {32'h446120db, 32'hc3c4f407} /* (18, 11, 1) {real, imag} */,
  {32'h44290298, 32'h00000000} /* (18, 11, 0) {real, imag} */,
  {32'hc446a058, 32'h4427788e} /* (18, 10, 31) {real, imag} */,
  {32'h43aa34ba, 32'hc2f113d8} /* (18, 10, 30) {real, imag} */,
  {32'h429723d1, 32'h42cf8aec} /* (18, 10, 29) {real, imag} */,
  {32'hc2cdebe5, 32'hc123efb0} /* (18, 10, 28) {real, imag} */,
  {32'h420b4872, 32'hc0de1470} /* (18, 10, 27) {real, imag} */,
  {32'hc2541c02, 32'h427d1c57} /* (18, 10, 26) {real, imag} */,
  {32'hc31965f3, 32'hc1e747ce} /* (18, 10, 25) {real, imag} */,
  {32'hc1864e39, 32'hc0ce6aa8} /* (18, 10, 24) {real, imag} */,
  {32'h406b8356, 32'hc1358dec} /* (18, 10, 23) {real, imag} */,
  {32'hc21a2cd8, 32'hc2c18e86} /* (18, 10, 22) {real, imag} */,
  {32'h41a1576b, 32'hc30b3cc6} /* (18, 10, 21) {real, imag} */,
  {32'h428bcd86, 32'hc166a75a} /* (18, 10, 20) {real, imag} */,
  {32'hc1e60a98, 32'h41f2d480} /* (18, 10, 19) {real, imag} */,
  {32'hc205254b, 32'hc24ec51a} /* (18, 10, 18) {real, imag} */,
  {32'h4288b779, 32'h424eb675} /* (18, 10, 17) {real, imag} */,
  {32'hbee51380, 32'h00000000} /* (18, 10, 16) {real, imag} */,
  {32'h4288b779, 32'hc24eb675} /* (18, 10, 15) {real, imag} */,
  {32'hc205254b, 32'h424ec51a} /* (18, 10, 14) {real, imag} */,
  {32'hc1e60a98, 32'hc1f2d480} /* (18, 10, 13) {real, imag} */,
  {32'h428bcd86, 32'h4166a75a} /* (18, 10, 12) {real, imag} */,
  {32'h41a1576b, 32'h430b3cc6} /* (18, 10, 11) {real, imag} */,
  {32'hc21a2cd8, 32'h42c18e86} /* (18, 10, 10) {real, imag} */,
  {32'h406b8356, 32'h41358dec} /* (18, 10, 9) {real, imag} */,
  {32'hc1864e39, 32'h40ce6aa8} /* (18, 10, 8) {real, imag} */,
  {32'hc31965f3, 32'h41e747ce} /* (18, 10, 7) {real, imag} */,
  {32'hc2541c02, 32'hc27d1c57} /* (18, 10, 6) {real, imag} */,
  {32'h420b4872, 32'h40de1470} /* (18, 10, 5) {real, imag} */,
  {32'hc2cdebe5, 32'h4123efb0} /* (18, 10, 4) {real, imag} */,
  {32'h429723d1, 32'hc2cf8aec} /* (18, 10, 3) {real, imag} */,
  {32'h43aa34ba, 32'h42f113d8} /* (18, 10, 2) {real, imag} */,
  {32'hc446a058, 32'hc427788e} /* (18, 10, 1) {real, imag} */,
  {32'hc438ba0c, 32'h00000000} /* (18, 10, 0) {real, imag} */,
  {32'hc5048248, 32'h44515b04} /* (18, 9, 31) {real, imag} */,
  {32'h445b67bd, 32'hc3688f44} /* (18, 9, 30) {real, imag} */,
  {32'hc231b0bc, 32'h4219e864} /* (18, 9, 29) {real, imag} */,
  {32'hc2715b12, 32'hc2095474} /* (18, 9, 28) {real, imag} */,
  {32'h427bacc4, 32'hc2898f10} /* (18, 9, 27) {real, imag} */,
  {32'h41a57740, 32'h42ce3b0f} /* (18, 9, 26) {real, imag} */,
  {32'hc2bd818e, 32'hc247d117} /* (18, 9, 25) {real, imag} */,
  {32'hc2b41698, 32'hc32063cc} /* (18, 9, 24) {real, imag} */,
  {32'h41f4591c, 32'hc28229f8} /* (18, 9, 23) {real, imag} */,
  {32'h40a22a78, 32'hc25073f8} /* (18, 9, 22) {real, imag} */,
  {32'h42a0433a, 32'hc2e62e66} /* (18, 9, 21) {real, imag} */,
  {32'h418d2fde, 32'hc2a5c062} /* (18, 9, 20) {real, imag} */,
  {32'hc18abaf0, 32'h427ad498} /* (18, 9, 19) {real, imag} */,
  {32'h41d4aeb3, 32'hc1de13b5} /* (18, 9, 18) {real, imag} */,
  {32'hc235f8a1, 32'hc1aa9d9c} /* (18, 9, 17) {real, imag} */,
  {32'hc2753a6a, 32'h00000000} /* (18, 9, 16) {real, imag} */,
  {32'hc235f8a1, 32'h41aa9d9c} /* (18, 9, 15) {real, imag} */,
  {32'h41d4aeb3, 32'h41de13b5} /* (18, 9, 14) {real, imag} */,
  {32'hc18abaf0, 32'hc27ad498} /* (18, 9, 13) {real, imag} */,
  {32'h418d2fde, 32'h42a5c062} /* (18, 9, 12) {real, imag} */,
  {32'h42a0433a, 32'h42e62e66} /* (18, 9, 11) {real, imag} */,
  {32'h40a22a78, 32'h425073f8} /* (18, 9, 10) {real, imag} */,
  {32'h41f4591c, 32'h428229f8} /* (18, 9, 9) {real, imag} */,
  {32'hc2b41698, 32'h432063cc} /* (18, 9, 8) {real, imag} */,
  {32'hc2bd818e, 32'h4247d117} /* (18, 9, 7) {real, imag} */,
  {32'h41a57740, 32'hc2ce3b0f} /* (18, 9, 6) {real, imag} */,
  {32'h427bacc4, 32'h42898f10} /* (18, 9, 5) {real, imag} */,
  {32'hc2715b12, 32'h42095474} /* (18, 9, 4) {real, imag} */,
  {32'hc231b0bc, 32'hc219e864} /* (18, 9, 3) {real, imag} */,
  {32'h445b67bd, 32'h43688f44} /* (18, 9, 2) {real, imag} */,
  {32'hc5048248, 32'hc4515b04} /* (18, 9, 1) {real, imag} */,
  {32'hc4e0f517, 32'h00000000} /* (18, 9, 0) {real, imag} */,
  {32'hc52d4c32, 32'h448c1332} /* (18, 8, 31) {real, imag} */,
  {32'h444ed6db, 32'hc3687928} /* (18, 8, 30) {real, imag} */,
  {32'h41f48742, 32'h42de3ac2} /* (18, 8, 29) {real, imag} */,
  {32'h422992a8, 32'h4114f858} /* (18, 8, 28) {real, imag} */,
  {32'h4317cce6, 32'hc2d9a173} /* (18, 8, 27) {real, imag} */,
  {32'h41e8441a, 32'h41ad4ea2} /* (18, 8, 26) {real, imag} */,
  {32'hc2a031d0, 32'h3f6ec3c0} /* (18, 8, 25) {real, imag} */,
  {32'h41e9c905, 32'hc2c223ff} /* (18, 8, 24) {real, imag} */,
  {32'h4081dca0, 32'h414bc873} /* (18, 8, 23) {real, imag} */,
  {32'hc2a537d8, 32'h42ed2487} /* (18, 8, 22) {real, imag} */,
  {32'h41057bc9, 32'h4288935a} /* (18, 8, 21) {real, imag} */,
  {32'hc1767bd4, 32'hc0d4f8c8} /* (18, 8, 20) {real, imag} */,
  {32'hc22a112c, 32'hc0bbc6e0} /* (18, 8, 19) {real, imag} */,
  {32'hc21d98e0, 32'hc2129e87} /* (18, 8, 18) {real, imag} */,
  {32'hc2a621b2, 32'h40c09366} /* (18, 8, 17) {real, imag} */,
  {32'hc1f5ffd1, 32'h00000000} /* (18, 8, 16) {real, imag} */,
  {32'hc2a621b2, 32'hc0c09366} /* (18, 8, 15) {real, imag} */,
  {32'hc21d98e0, 32'h42129e87} /* (18, 8, 14) {real, imag} */,
  {32'hc22a112c, 32'h40bbc6e0} /* (18, 8, 13) {real, imag} */,
  {32'hc1767bd4, 32'h40d4f8c8} /* (18, 8, 12) {real, imag} */,
  {32'h41057bc9, 32'hc288935a} /* (18, 8, 11) {real, imag} */,
  {32'hc2a537d8, 32'hc2ed2487} /* (18, 8, 10) {real, imag} */,
  {32'h4081dca0, 32'hc14bc873} /* (18, 8, 9) {real, imag} */,
  {32'h41e9c905, 32'h42c223ff} /* (18, 8, 8) {real, imag} */,
  {32'hc2a031d0, 32'hbf6ec3c0} /* (18, 8, 7) {real, imag} */,
  {32'h41e8441a, 32'hc1ad4ea2} /* (18, 8, 6) {real, imag} */,
  {32'h4317cce6, 32'h42d9a173} /* (18, 8, 5) {real, imag} */,
  {32'h422992a8, 32'hc114f858} /* (18, 8, 4) {real, imag} */,
  {32'h41f48742, 32'hc2de3ac2} /* (18, 8, 3) {real, imag} */,
  {32'h444ed6db, 32'h43687928} /* (18, 8, 2) {real, imag} */,
  {32'hc52d4c32, 32'hc48c1332} /* (18, 8, 1) {real, imag} */,
  {32'hc51d1008, 32'h00000000} /* (18, 8, 0) {real, imag} */,
  {32'hc5404dca, 32'h44b85ac2} /* (18, 7, 31) {real, imag} */,
  {32'h447bf831, 32'hc3bb8560} /* (18, 7, 30) {real, imag} */,
  {32'hc1d7bd22, 32'h415377f4} /* (18, 7, 29) {real, imag} */,
  {32'hc2f96e40, 32'h42a873da} /* (18, 7, 28) {real, imag} */,
  {32'h41c94628, 32'hc2e6903c} /* (18, 7, 27) {real, imag} */,
  {32'hc1f6a238, 32'h43024004} /* (18, 7, 26) {real, imag} */,
  {32'hc22548d0, 32'hc1fc75ec} /* (18, 7, 25) {real, imag} */,
  {32'h4222f349, 32'hc389482b} /* (18, 7, 24) {real, imag} */,
  {32'h418a9529, 32'h42bdc151} /* (18, 7, 23) {real, imag} */,
  {32'hc1d0a056, 32'h42070a78} /* (18, 7, 22) {real, imag} */,
  {32'h4283c6ae, 32'hc24a9d5a} /* (18, 7, 21) {real, imag} */,
  {32'hc15fcd0c, 32'hc26eb741} /* (18, 7, 20) {real, imag} */,
  {32'h427fdad7, 32'hc1771958} /* (18, 7, 19) {real, imag} */,
  {32'hc0385620, 32'hc2b83e99} /* (18, 7, 18) {real, imag} */,
  {32'h41d79c35, 32'h43048408} /* (18, 7, 17) {real, imag} */,
  {32'h41e96406, 32'h00000000} /* (18, 7, 16) {real, imag} */,
  {32'h41d79c35, 32'hc3048408} /* (18, 7, 15) {real, imag} */,
  {32'hc0385620, 32'h42b83e99} /* (18, 7, 14) {real, imag} */,
  {32'h427fdad7, 32'h41771958} /* (18, 7, 13) {real, imag} */,
  {32'hc15fcd0c, 32'h426eb741} /* (18, 7, 12) {real, imag} */,
  {32'h4283c6ae, 32'h424a9d5a} /* (18, 7, 11) {real, imag} */,
  {32'hc1d0a056, 32'hc2070a78} /* (18, 7, 10) {real, imag} */,
  {32'h418a9529, 32'hc2bdc151} /* (18, 7, 9) {real, imag} */,
  {32'h4222f349, 32'h4389482b} /* (18, 7, 8) {real, imag} */,
  {32'hc22548d0, 32'h41fc75ec} /* (18, 7, 7) {real, imag} */,
  {32'hc1f6a238, 32'hc3024004} /* (18, 7, 6) {real, imag} */,
  {32'h41c94628, 32'h42e6903c} /* (18, 7, 5) {real, imag} */,
  {32'hc2f96e40, 32'hc2a873da} /* (18, 7, 4) {real, imag} */,
  {32'hc1d7bd22, 32'hc15377f4} /* (18, 7, 3) {real, imag} */,
  {32'h447bf831, 32'h43bb8560} /* (18, 7, 2) {real, imag} */,
  {32'hc5404dca, 32'hc4b85ac2} /* (18, 7, 1) {real, imag} */,
  {32'hc53b12ee, 32'h00000000} /* (18, 7, 0) {real, imag} */,
  {32'hc546c8a0, 32'h44eaece2} /* (18, 6, 31) {real, imag} */,
  {32'h4436498a, 32'hc433b64e} /* (18, 6, 30) {real, imag} */,
  {32'hc2dce935, 32'hc333bb16} /* (18, 6, 29) {real, imag} */,
  {32'hc281e822, 32'h429ccd1d} /* (18, 6, 28) {real, imag} */,
  {32'h433fa193, 32'hc1d274da} /* (18, 6, 27) {real, imag} */,
  {32'h4294aea1, 32'h42defaaa} /* (18, 6, 26) {real, imag} */,
  {32'h4340601c, 32'h4204190e} /* (18, 6, 25) {real, imag} */,
  {32'h42cb0b56, 32'hc31e402c} /* (18, 6, 24) {real, imag} */,
  {32'hc0bfed22, 32'hc184956e} /* (18, 6, 23) {real, imag} */,
  {32'h4127e574, 32'h41210414} /* (18, 6, 22) {real, imag} */,
  {32'h41b24219, 32'h41840349} /* (18, 6, 21) {real, imag} */,
  {32'hc2ed4122, 32'h4230e704} /* (18, 6, 20) {real, imag} */,
  {32'h41c0e910, 32'hc219b276} /* (18, 6, 19) {real, imag} */,
  {32'hc2c997a9, 32'h412a2be6} /* (18, 6, 18) {real, imag} */,
  {32'hc117b894, 32'h4216e531} /* (18, 6, 17) {real, imag} */,
  {32'hc08221f8, 32'h00000000} /* (18, 6, 16) {real, imag} */,
  {32'hc117b894, 32'hc216e531} /* (18, 6, 15) {real, imag} */,
  {32'hc2c997a9, 32'hc12a2be6} /* (18, 6, 14) {real, imag} */,
  {32'h41c0e910, 32'h4219b276} /* (18, 6, 13) {real, imag} */,
  {32'hc2ed4122, 32'hc230e704} /* (18, 6, 12) {real, imag} */,
  {32'h41b24219, 32'hc1840349} /* (18, 6, 11) {real, imag} */,
  {32'h4127e574, 32'hc1210414} /* (18, 6, 10) {real, imag} */,
  {32'hc0bfed22, 32'h4184956e} /* (18, 6, 9) {real, imag} */,
  {32'h42cb0b56, 32'h431e402c} /* (18, 6, 8) {real, imag} */,
  {32'h4340601c, 32'hc204190e} /* (18, 6, 7) {real, imag} */,
  {32'h4294aea1, 32'hc2defaaa} /* (18, 6, 6) {real, imag} */,
  {32'h433fa193, 32'h41d274da} /* (18, 6, 5) {real, imag} */,
  {32'hc281e822, 32'hc29ccd1d} /* (18, 6, 4) {real, imag} */,
  {32'hc2dce935, 32'h4333bb16} /* (18, 6, 3) {real, imag} */,
  {32'h4436498a, 32'h4433b64e} /* (18, 6, 2) {real, imag} */,
  {32'hc546c8a0, 32'hc4eaece2} /* (18, 6, 1) {real, imag} */,
  {32'hc54c8518, 32'h00000000} /* (18, 6, 0) {real, imag} */,
  {32'hc52ee7e7, 32'h45173a92} /* (18, 5, 31) {real, imag} */,
  {32'h435086e8, 32'hc4595ada} /* (18, 5, 30) {real, imag} */,
  {32'hc08e2df4, 32'hc2926023} /* (18, 5, 29) {real, imag} */,
  {32'h428a676c, 32'hc240c7e2} /* (18, 5, 28) {real, imag} */,
  {32'h431fd6d2, 32'h421de413} /* (18, 5, 27) {real, imag} */,
  {32'h4308d01c, 32'hc23c0b7c} /* (18, 5, 26) {real, imag} */,
  {32'hc0a80044, 32'hc1e3cab4} /* (18, 5, 25) {real, imag} */,
  {32'h425b15ac, 32'h41ea8f4a} /* (18, 5, 24) {real, imag} */,
  {32'hc209b546, 32'hc2d49ef2} /* (18, 5, 23) {real, imag} */,
  {32'hc2c2a4e2, 32'h4280ca76} /* (18, 5, 22) {real, imag} */,
  {32'hc248a00d, 32'h42d43f08} /* (18, 5, 21) {real, imag} */,
  {32'h426f95a3, 32'hc2bbad7e} /* (18, 5, 20) {real, imag} */,
  {32'h41b03361, 32'h41bae7f8} /* (18, 5, 19) {real, imag} */,
  {32'h3fbb8490, 32'h4261cbc4} /* (18, 5, 18) {real, imag} */,
  {32'h4230e7ec, 32'h413fa02e} /* (18, 5, 17) {real, imag} */,
  {32'h41155fc5, 32'h00000000} /* (18, 5, 16) {real, imag} */,
  {32'h4230e7ec, 32'hc13fa02e} /* (18, 5, 15) {real, imag} */,
  {32'h3fbb8490, 32'hc261cbc4} /* (18, 5, 14) {real, imag} */,
  {32'h41b03361, 32'hc1bae7f8} /* (18, 5, 13) {real, imag} */,
  {32'h426f95a3, 32'h42bbad7e} /* (18, 5, 12) {real, imag} */,
  {32'hc248a00d, 32'hc2d43f08} /* (18, 5, 11) {real, imag} */,
  {32'hc2c2a4e2, 32'hc280ca76} /* (18, 5, 10) {real, imag} */,
  {32'hc209b546, 32'h42d49ef2} /* (18, 5, 9) {real, imag} */,
  {32'h425b15ac, 32'hc1ea8f4a} /* (18, 5, 8) {real, imag} */,
  {32'hc0a80044, 32'h41e3cab4} /* (18, 5, 7) {real, imag} */,
  {32'h4308d01c, 32'h423c0b7c} /* (18, 5, 6) {real, imag} */,
  {32'h431fd6d2, 32'hc21de413} /* (18, 5, 5) {real, imag} */,
  {32'h428a676c, 32'h4240c7e2} /* (18, 5, 4) {real, imag} */,
  {32'hc08e2df4, 32'h42926023} /* (18, 5, 3) {real, imag} */,
  {32'h435086e8, 32'h44595ada} /* (18, 5, 2) {real, imag} */,
  {32'hc52ee7e7, 32'hc5173a92} /* (18, 5, 1) {real, imag} */,
  {32'hc560977a, 32'h00000000} /* (18, 5, 0) {real, imag} */,
  {32'hc51de71f, 32'h453533e8} /* (18, 4, 31) {real, imag} */,
  {32'hc3560e84, 32'hc4885a4d} /* (18, 4, 30) {real, imag} */,
  {32'h426dde58, 32'hc214c1cc} /* (18, 4, 29) {real, imag} */,
  {32'h43729189, 32'h41ee158e} /* (18, 4, 28) {real, imag} */,
  {32'h434b426d, 32'h42f4ebb6} /* (18, 4, 27) {real, imag} */,
  {32'h4306917f, 32'h4127a93e} /* (18, 4, 26) {real, imag} */,
  {32'hc24b44f0, 32'h4222ab2c} /* (18, 4, 25) {real, imag} */,
  {32'hc1b14fbd, 32'hc2b0cec7} /* (18, 4, 24) {real, imag} */,
  {32'hc1596700, 32'hc2977a38} /* (18, 4, 23) {real, imag} */,
  {32'hc0c0f968, 32'hc2baee18} /* (18, 4, 22) {real, imag} */,
  {32'hc1930610, 32'h41273c84} /* (18, 4, 21) {real, imag} */,
  {32'hc1d4da34, 32'hc1a2df66} /* (18, 4, 20) {real, imag} */,
  {32'h41eef610, 32'h40be0080} /* (18, 4, 19) {real, imag} */,
  {32'h4280f372, 32'hc29acf57} /* (18, 4, 18) {real, imag} */,
  {32'hc0d976cc, 32'h427040b6} /* (18, 4, 17) {real, imag} */,
  {32'h426765fb, 32'h00000000} /* (18, 4, 16) {real, imag} */,
  {32'hc0d976cc, 32'hc27040b6} /* (18, 4, 15) {real, imag} */,
  {32'h4280f372, 32'h429acf57} /* (18, 4, 14) {real, imag} */,
  {32'h41eef610, 32'hc0be0080} /* (18, 4, 13) {real, imag} */,
  {32'hc1d4da34, 32'h41a2df66} /* (18, 4, 12) {real, imag} */,
  {32'hc1930610, 32'hc1273c84} /* (18, 4, 11) {real, imag} */,
  {32'hc0c0f968, 32'h42baee18} /* (18, 4, 10) {real, imag} */,
  {32'hc1596700, 32'h42977a38} /* (18, 4, 9) {real, imag} */,
  {32'hc1b14fbd, 32'h42b0cec7} /* (18, 4, 8) {real, imag} */,
  {32'hc24b44f0, 32'hc222ab2c} /* (18, 4, 7) {real, imag} */,
  {32'h4306917f, 32'hc127a93e} /* (18, 4, 6) {real, imag} */,
  {32'h434b426d, 32'hc2f4ebb6} /* (18, 4, 5) {real, imag} */,
  {32'h43729189, 32'hc1ee158e} /* (18, 4, 4) {real, imag} */,
  {32'h426dde58, 32'h4214c1cc} /* (18, 4, 3) {real, imag} */,
  {32'hc3560e84, 32'h44885a4d} /* (18, 4, 2) {real, imag} */,
  {32'hc51de71f, 32'hc53533e8} /* (18, 4, 1) {real, imag} */,
  {32'hc567928d, 32'h00000000} /* (18, 4, 0) {real, imag} */,
  {32'hc517395a, 32'h453c9420} /* (18, 3, 31) {real, imag} */,
  {32'hc3b1b311, 32'hc4941cf2} /* (18, 3, 30) {real, imag} */,
  {32'h41c9949c, 32'hc22f5a0b} /* (18, 3, 29) {real, imag} */,
  {32'h42852b4b, 32'hc308bd40} /* (18, 3, 28) {real, imag} */,
  {32'h4381621d, 32'h42e9697b} /* (18, 3, 27) {real, imag} */,
  {32'h4192e878, 32'hc23198bc} /* (18, 3, 26) {real, imag} */,
  {32'hc142c1b0, 32'h42c0416e} /* (18, 3, 25) {real, imag} */,
  {32'h4274532c, 32'hc2143dc6} /* (18, 3, 24) {real, imag} */,
  {32'hc2106a19, 32'hc2785d41} /* (18, 3, 23) {real, imag} */,
  {32'hc1b67196, 32'hc2968b61} /* (18, 3, 22) {real, imag} */,
  {32'h43039d34, 32'h403748b0} /* (18, 3, 21) {real, imag} */,
  {32'h40f60b58, 32'hc1eedd63} /* (18, 3, 20) {real, imag} */,
  {32'hc11c461a, 32'hc1af324f} /* (18, 3, 19) {real, imag} */,
  {32'h40fcbc9b, 32'h41a720ca} /* (18, 3, 18) {real, imag} */,
  {32'h3f246940, 32'h4172a49b} /* (18, 3, 17) {real, imag} */,
  {32'h4238b576, 32'h00000000} /* (18, 3, 16) {real, imag} */,
  {32'h3f246940, 32'hc172a49b} /* (18, 3, 15) {real, imag} */,
  {32'h40fcbc9b, 32'hc1a720ca} /* (18, 3, 14) {real, imag} */,
  {32'hc11c461a, 32'h41af324f} /* (18, 3, 13) {real, imag} */,
  {32'h40f60b58, 32'h41eedd63} /* (18, 3, 12) {real, imag} */,
  {32'h43039d34, 32'hc03748b0} /* (18, 3, 11) {real, imag} */,
  {32'hc1b67196, 32'h42968b61} /* (18, 3, 10) {real, imag} */,
  {32'hc2106a19, 32'h42785d41} /* (18, 3, 9) {real, imag} */,
  {32'h4274532c, 32'h42143dc6} /* (18, 3, 8) {real, imag} */,
  {32'hc142c1b0, 32'hc2c0416e} /* (18, 3, 7) {real, imag} */,
  {32'h4192e878, 32'h423198bc} /* (18, 3, 6) {real, imag} */,
  {32'h4381621d, 32'hc2e9697b} /* (18, 3, 5) {real, imag} */,
  {32'h42852b4b, 32'h4308bd40} /* (18, 3, 4) {real, imag} */,
  {32'h41c9949c, 32'h422f5a0b} /* (18, 3, 3) {real, imag} */,
  {32'hc3b1b311, 32'h44941cf2} /* (18, 3, 2) {real, imag} */,
  {32'hc517395a, 32'hc53c9420} /* (18, 3, 1) {real, imag} */,
  {32'hc5655107, 32'h00000000} /* (18, 3, 0) {real, imag} */,
  {32'hc5133630, 32'h45398ede} /* (18, 2, 31) {real, imag} */,
  {32'hc3d4f5b7, 32'hc48a9220} /* (18, 2, 30) {real, imag} */,
  {32'h42f86db3, 32'hc1c31cd8} /* (18, 2, 29) {real, imag} */,
  {32'h42d3bbc3, 32'hc383f6ee} /* (18, 2, 28) {real, imag} */,
  {32'h432253d8, 32'h432a7d92} /* (18, 2, 27) {real, imag} */,
  {32'hc00304a0, 32'hc1f2264a} /* (18, 2, 26) {real, imag} */,
  {32'hc26aa5da, 32'h413121d8} /* (18, 2, 25) {real, imag} */,
  {32'h425ee9fe, 32'h3f2e1b40} /* (18, 2, 24) {real, imag} */,
  {32'h42c1df95, 32'hc2c5561e} /* (18, 2, 23) {real, imag} */,
  {32'h4267415c, 32'hc1f9a1b3} /* (18, 2, 22) {real, imag} */,
  {32'h42d13a3c, 32'h40fc1d00} /* (18, 2, 21) {real, imag} */,
  {32'hc11a2532, 32'hc29b39b0} /* (18, 2, 20) {real, imag} */,
  {32'h427eda64, 32'h41ce66be} /* (18, 2, 19) {real, imag} */,
  {32'hc2fed610, 32'hc22ce3ad} /* (18, 2, 18) {real, imag} */,
  {32'h424cd323, 32'hc1614196} /* (18, 2, 17) {real, imag} */,
  {32'h41b8a754, 32'h00000000} /* (18, 2, 16) {real, imag} */,
  {32'h424cd323, 32'h41614196} /* (18, 2, 15) {real, imag} */,
  {32'hc2fed610, 32'h422ce3ad} /* (18, 2, 14) {real, imag} */,
  {32'h427eda64, 32'hc1ce66be} /* (18, 2, 13) {real, imag} */,
  {32'hc11a2532, 32'h429b39b0} /* (18, 2, 12) {real, imag} */,
  {32'h42d13a3c, 32'hc0fc1d00} /* (18, 2, 11) {real, imag} */,
  {32'h4267415c, 32'h41f9a1b3} /* (18, 2, 10) {real, imag} */,
  {32'h42c1df95, 32'h42c5561e} /* (18, 2, 9) {real, imag} */,
  {32'h425ee9fe, 32'hbf2e1b40} /* (18, 2, 8) {real, imag} */,
  {32'hc26aa5da, 32'hc13121d8} /* (18, 2, 7) {real, imag} */,
  {32'hc00304a0, 32'h41f2264a} /* (18, 2, 6) {real, imag} */,
  {32'h432253d8, 32'hc32a7d92} /* (18, 2, 5) {real, imag} */,
  {32'h42d3bbc3, 32'h4383f6ee} /* (18, 2, 4) {real, imag} */,
  {32'h42f86db3, 32'h41c31cd8} /* (18, 2, 3) {real, imag} */,
  {32'hc3d4f5b7, 32'h448a9220} /* (18, 2, 2) {real, imag} */,
  {32'hc5133630, 32'hc5398ede} /* (18, 2, 1) {real, imag} */,
  {32'hc5727bbf, 32'h00000000} /* (18, 2, 0) {real, imag} */,
  {32'hc51bec4f, 32'h452afb01} /* (18, 1, 31) {real, imag} */,
  {32'hc396a812, 32'hc47df188} /* (18, 1, 30) {real, imag} */,
  {32'h43081d22, 32'h42affa3a} /* (18, 1, 29) {real, imag} */,
  {32'h41b27aa9, 32'hc391f218} /* (18, 1, 28) {real, imag} */,
  {32'h431e144a, 32'h430d1c63} /* (18, 1, 27) {real, imag} */,
  {32'h43192cc0, 32'hc2806d78} /* (18, 1, 26) {real, imag} */,
  {32'h41c137f6, 32'hc1158276} /* (18, 1, 25) {real, imag} */,
  {32'h42d2e7b4, 32'hc1ae8fe4} /* (18, 1, 24) {real, imag} */,
  {32'h41d8c1ad, 32'h418737a7} /* (18, 1, 23) {real, imag} */,
  {32'h4182358f, 32'h41f48784} /* (18, 1, 22) {real, imag} */,
  {32'h416ca704, 32'hc0a2a7b8} /* (18, 1, 21) {real, imag} */,
  {32'h412ad9b2, 32'h41f2a36a} /* (18, 1, 20) {real, imag} */,
  {32'hc1d81014, 32'h424437d8} /* (18, 1, 19) {real, imag} */,
  {32'hc20236b5, 32'h4055d190} /* (18, 1, 18) {real, imag} */,
  {32'h41d364e1, 32'h41e5a60d} /* (18, 1, 17) {real, imag} */,
  {32'h40f0ad5c, 32'h00000000} /* (18, 1, 16) {real, imag} */,
  {32'h41d364e1, 32'hc1e5a60d} /* (18, 1, 15) {real, imag} */,
  {32'hc20236b5, 32'hc055d190} /* (18, 1, 14) {real, imag} */,
  {32'hc1d81014, 32'hc24437d8} /* (18, 1, 13) {real, imag} */,
  {32'h412ad9b2, 32'hc1f2a36a} /* (18, 1, 12) {real, imag} */,
  {32'h416ca704, 32'h40a2a7b8} /* (18, 1, 11) {real, imag} */,
  {32'h4182358f, 32'hc1f48784} /* (18, 1, 10) {real, imag} */,
  {32'h41d8c1ad, 32'hc18737a7} /* (18, 1, 9) {real, imag} */,
  {32'h42d2e7b4, 32'h41ae8fe4} /* (18, 1, 8) {real, imag} */,
  {32'h41c137f6, 32'h41158276} /* (18, 1, 7) {real, imag} */,
  {32'h43192cc0, 32'h42806d78} /* (18, 1, 6) {real, imag} */,
  {32'h431e144a, 32'hc30d1c63} /* (18, 1, 5) {real, imag} */,
  {32'h41b27aa9, 32'h4391f218} /* (18, 1, 4) {real, imag} */,
  {32'h43081d22, 32'hc2affa3a} /* (18, 1, 3) {real, imag} */,
  {32'hc396a812, 32'h447df188} /* (18, 1, 2) {real, imag} */,
  {32'hc51bec4f, 32'hc52afb01} /* (18, 1, 1) {real, imag} */,
  {32'hc5794a06, 32'h00000000} /* (18, 1, 0) {real, imag} */,
  {32'hc52a71c4, 32'h450b0ae4} /* (18, 0, 31) {real, imag} */,
  {32'h41a56ae0, 32'hc434e6a2} /* (18, 0, 30) {real, imag} */,
  {32'h413bdd10, 32'h42676d34} /* (18, 0, 29) {real, imag} */,
  {32'hc0dd8840, 32'hc318d88c} /* (18, 0, 28) {real, imag} */,
  {32'h42ac61fa, 32'hc176d090} /* (18, 0, 27) {real, imag} */,
  {32'hbfbc1230, 32'hc21d74e1} /* (18, 0, 26) {real, imag} */,
  {32'h41931ddb, 32'h41c4f868} /* (18, 0, 25) {real, imag} */,
  {32'h426fdc78, 32'hc2b14b32} /* (18, 0, 24) {real, imag} */,
  {32'hc074823c, 32'h42792196} /* (18, 0, 23) {real, imag} */,
  {32'h4188c5a7, 32'hc2466b32} /* (18, 0, 22) {real, imag} */,
  {32'hc191cf74, 32'hc208caff} /* (18, 0, 21) {real, imag} */,
  {32'h427fb774, 32'hc1d1acbd} /* (18, 0, 20) {real, imag} */,
  {32'h428e445b, 32'h4191eb1c} /* (18, 0, 19) {real, imag} */,
  {32'h42189fe5, 32'h41ee0e38} /* (18, 0, 18) {real, imag} */,
  {32'h41847792, 32'hc0c50b92} /* (18, 0, 17) {real, imag} */,
  {32'hc1a83c14, 32'h00000000} /* (18, 0, 16) {real, imag} */,
  {32'h41847792, 32'h40c50b92} /* (18, 0, 15) {real, imag} */,
  {32'h42189fe5, 32'hc1ee0e38} /* (18, 0, 14) {real, imag} */,
  {32'h428e445b, 32'hc191eb1c} /* (18, 0, 13) {real, imag} */,
  {32'h427fb774, 32'h41d1acbd} /* (18, 0, 12) {real, imag} */,
  {32'hc191cf74, 32'h4208caff} /* (18, 0, 11) {real, imag} */,
  {32'h4188c5a7, 32'h42466b32} /* (18, 0, 10) {real, imag} */,
  {32'hc074823c, 32'hc2792196} /* (18, 0, 9) {real, imag} */,
  {32'h426fdc78, 32'h42b14b32} /* (18, 0, 8) {real, imag} */,
  {32'h41931ddb, 32'hc1c4f868} /* (18, 0, 7) {real, imag} */,
  {32'hbfbc1230, 32'h421d74e1} /* (18, 0, 6) {real, imag} */,
  {32'h42ac61fa, 32'h4176d090} /* (18, 0, 5) {real, imag} */,
  {32'hc0dd8840, 32'h4318d88c} /* (18, 0, 4) {real, imag} */,
  {32'h413bdd10, 32'hc2676d34} /* (18, 0, 3) {real, imag} */,
  {32'h41a56ae0, 32'h4434e6a2} /* (18, 0, 2) {real, imag} */,
  {32'hc52a71c4, 32'hc50b0ae4} /* (18, 0, 1) {real, imag} */,
  {32'hc567dd84, 32'h00000000} /* (18, 0, 0) {real, imag} */,
  {32'hc507eb98, 32'h448ad737} /* (17, 31, 31) {real, imag} */,
  {32'h43e92877, 32'hc3f23056} /* (17, 31, 30) {real, imag} */,
  {32'h4246adae, 32'h421737b6} /* (17, 31, 29) {real, imag} */,
  {32'hc2041f2a, 32'h418e6fd0} /* (17, 31, 28) {real, imag} */,
  {32'h4278ecf2, 32'hc2385544} /* (17, 31, 27) {real, imag} */,
  {32'h425eb6eb, 32'h40734710} /* (17, 31, 26) {real, imag} */,
  {32'h41880512, 32'h40d38388} /* (17, 31, 25) {real, imag} */,
  {32'hc1f85a89, 32'hc2511308} /* (17, 31, 24) {real, imag} */,
  {32'hbfa77fd0, 32'h418912d2} /* (17, 31, 23) {real, imag} */,
  {32'h413108f0, 32'h41e23736} /* (17, 31, 22) {real, imag} */,
  {32'h42827b4c, 32'hc26b62df} /* (17, 31, 21) {real, imag} */,
  {32'hc10e136c, 32'h40927b60} /* (17, 31, 20) {real, imag} */,
  {32'h41f8a8a5, 32'h416c3ff7} /* (17, 31, 19) {real, imag} */,
  {32'hc2957e63, 32'hc0b5ba78} /* (17, 31, 18) {real, imag} */,
  {32'h4234a4f0, 32'hc15a37e2} /* (17, 31, 17) {real, imag} */,
  {32'hc08674ac, 32'h00000000} /* (17, 31, 16) {real, imag} */,
  {32'h4234a4f0, 32'h415a37e2} /* (17, 31, 15) {real, imag} */,
  {32'hc2957e63, 32'h40b5ba78} /* (17, 31, 14) {real, imag} */,
  {32'h41f8a8a5, 32'hc16c3ff7} /* (17, 31, 13) {real, imag} */,
  {32'hc10e136c, 32'hc0927b60} /* (17, 31, 12) {real, imag} */,
  {32'h42827b4c, 32'h426b62df} /* (17, 31, 11) {real, imag} */,
  {32'h413108f0, 32'hc1e23736} /* (17, 31, 10) {real, imag} */,
  {32'hbfa77fd0, 32'hc18912d2} /* (17, 31, 9) {real, imag} */,
  {32'hc1f85a89, 32'h42511308} /* (17, 31, 8) {real, imag} */,
  {32'h41880512, 32'hc0d38388} /* (17, 31, 7) {real, imag} */,
  {32'h425eb6eb, 32'hc0734710} /* (17, 31, 6) {real, imag} */,
  {32'h4278ecf2, 32'h42385544} /* (17, 31, 5) {real, imag} */,
  {32'hc2041f2a, 32'hc18e6fd0} /* (17, 31, 4) {real, imag} */,
  {32'h4246adae, 32'hc21737b6} /* (17, 31, 3) {real, imag} */,
  {32'h43e92877, 32'h43f23056} /* (17, 31, 2) {real, imag} */,
  {32'hc507eb98, 32'hc48ad737} /* (17, 31, 1) {real, imag} */,
  {32'hc52253aa, 32'h00000000} /* (17, 31, 0) {real, imag} */,
  {32'hc52d42b2, 32'h4441df68} /* (17, 30, 31) {real, imag} */,
  {32'h444b3d3f, 32'hc3d27684} /* (17, 30, 30) {real, imag} */,
  {32'h41bfac50, 32'h429cb4a4} /* (17, 30, 29) {real, imag} */,
  {32'hc2d09e50, 32'h42dc7b26} /* (17, 30, 28) {real, imag} */,
  {32'h4381cff2, 32'hc225bc6c} /* (17, 30, 27) {real, imag} */,
  {32'h4286666c, 32'hc2a58990} /* (17, 30, 26) {real, imag} */,
  {32'h422b689c, 32'hc1968a88} /* (17, 30, 25) {real, imag} */,
  {32'h429ef7b0, 32'hc3065407} /* (17, 30, 24) {real, imag} */,
  {32'hc283e182, 32'h4299d4ac} /* (17, 30, 23) {real, imag} */,
  {32'h422673df, 32'h4225b215} /* (17, 30, 22) {real, imag} */,
  {32'h422baea4, 32'hc1b4f328} /* (17, 30, 21) {real, imag} */,
  {32'hc1336ddc, 32'h425c08f4} /* (17, 30, 20) {real, imag} */,
  {32'h41534bec, 32'h41f65f81} /* (17, 30, 19) {real, imag} */,
  {32'hc1db8596, 32'hc0a7d0cc} /* (17, 30, 18) {real, imag} */,
  {32'hc14cfe44, 32'h4208682c} /* (17, 30, 17) {real, imag} */,
  {32'hc13fc278, 32'h00000000} /* (17, 30, 16) {real, imag} */,
  {32'hc14cfe44, 32'hc208682c} /* (17, 30, 15) {real, imag} */,
  {32'hc1db8596, 32'h40a7d0cc} /* (17, 30, 14) {real, imag} */,
  {32'h41534bec, 32'hc1f65f81} /* (17, 30, 13) {real, imag} */,
  {32'hc1336ddc, 32'hc25c08f4} /* (17, 30, 12) {real, imag} */,
  {32'h422baea4, 32'h41b4f328} /* (17, 30, 11) {real, imag} */,
  {32'h422673df, 32'hc225b215} /* (17, 30, 10) {real, imag} */,
  {32'hc283e182, 32'hc299d4ac} /* (17, 30, 9) {real, imag} */,
  {32'h429ef7b0, 32'h43065407} /* (17, 30, 8) {real, imag} */,
  {32'h422b689c, 32'h41968a88} /* (17, 30, 7) {real, imag} */,
  {32'h4286666c, 32'h42a58990} /* (17, 30, 6) {real, imag} */,
  {32'h4381cff2, 32'h4225bc6c} /* (17, 30, 5) {real, imag} */,
  {32'hc2d09e50, 32'hc2dc7b26} /* (17, 30, 4) {real, imag} */,
  {32'h41bfac50, 32'hc29cb4a4} /* (17, 30, 3) {real, imag} */,
  {32'h444b3d3f, 32'h43d27684} /* (17, 30, 2) {real, imag} */,
  {32'hc52d42b2, 32'hc441df68} /* (17, 30, 1) {real, imag} */,
  {32'hc52e1a99, 32'h00000000} /* (17, 30, 0) {real, imag} */,
  {32'hc5442b02, 32'h4427b7e8} /* (17, 29, 31) {real, imag} */,
  {32'h44833d6f, 32'hc3ad2b6b} /* (17, 29, 30) {real, imag} */,
  {32'hc2a52ede, 32'h42c850a8} /* (17, 29, 29) {real, imag} */,
  {32'hc33ce1c0, 32'h42e30058} /* (17, 29, 28) {real, imag} */,
  {32'h434f0498, 32'hc21492f0} /* (17, 29, 27) {real, imag} */,
  {32'h42fcf2ca, 32'hc0d47620} /* (17, 29, 26) {real, imag} */,
  {32'hc260a7f7, 32'h3fbc9980} /* (17, 29, 25) {real, imag} */,
  {32'h42328b52, 32'hc1acb088} /* (17, 29, 24) {real, imag} */,
  {32'hc2e5019e, 32'hc2acf9b8} /* (17, 29, 23) {real, imag} */,
  {32'h42bbea76, 32'h42066546} /* (17, 29, 22) {real, imag} */,
  {32'hc19fc100, 32'hc0c91cf0} /* (17, 29, 21) {real, imag} */,
  {32'hc2cd4bdc, 32'h3f95cb98} /* (17, 29, 20) {real, imag} */,
  {32'h4106b8a9, 32'h420bdc08} /* (17, 29, 19) {real, imag} */,
  {32'hc10e3b44, 32'hc1c0fd4a} /* (17, 29, 18) {real, imag} */,
  {32'hc1b8262d, 32'h41a6156a} /* (17, 29, 17) {real, imag} */,
  {32'hc2de41b4, 32'h00000000} /* (17, 29, 16) {real, imag} */,
  {32'hc1b8262d, 32'hc1a6156a} /* (17, 29, 15) {real, imag} */,
  {32'hc10e3b44, 32'h41c0fd4a} /* (17, 29, 14) {real, imag} */,
  {32'h4106b8a9, 32'hc20bdc08} /* (17, 29, 13) {real, imag} */,
  {32'hc2cd4bdc, 32'hbf95cb98} /* (17, 29, 12) {real, imag} */,
  {32'hc19fc100, 32'h40c91cf0} /* (17, 29, 11) {real, imag} */,
  {32'h42bbea76, 32'hc2066546} /* (17, 29, 10) {real, imag} */,
  {32'hc2e5019e, 32'h42acf9b8} /* (17, 29, 9) {real, imag} */,
  {32'h42328b52, 32'h41acb088} /* (17, 29, 8) {real, imag} */,
  {32'hc260a7f7, 32'hbfbc9980} /* (17, 29, 7) {real, imag} */,
  {32'h42fcf2ca, 32'h40d47620} /* (17, 29, 6) {real, imag} */,
  {32'h434f0498, 32'h421492f0} /* (17, 29, 5) {real, imag} */,
  {32'hc33ce1c0, 32'hc2e30058} /* (17, 29, 4) {real, imag} */,
  {32'hc2a52ede, 32'hc2c850a8} /* (17, 29, 3) {real, imag} */,
  {32'h44833d6f, 32'h43ad2b6b} /* (17, 29, 2) {real, imag} */,
  {32'hc5442b02, 32'hc427b7e8} /* (17, 29, 1) {real, imag} */,
  {32'hc53331de, 32'h00000000} /* (17, 29, 0) {real, imag} */,
  {32'hc549b455, 32'h4413a116} /* (17, 28, 31) {real, imag} */,
  {32'h4482c906, 32'hc3cf5d1a} /* (17, 28, 30) {real, imag} */,
  {32'hc160cd28, 32'hc1a8bce7} /* (17, 28, 29) {real, imag} */,
  {32'hc3261405, 32'h426b8e36} /* (17, 28, 28) {real, imag} */,
  {32'h430b90b6, 32'hc25211ec} /* (17, 28, 27) {real, imag} */,
  {32'h430ab31d, 32'h4113387a} /* (17, 28, 26) {real, imag} */,
  {32'hc0fe3508, 32'hc215e397} /* (17, 28, 25) {real, imag} */,
  {32'h41bbcf82, 32'hc1c6b734} /* (17, 28, 24) {real, imag} */,
  {32'h42820c4a, 32'h41fb97e1} /* (17, 28, 23) {real, imag} */,
  {32'h4185858f, 32'h41048348} /* (17, 28, 22) {real, imag} */,
  {32'h42592726, 32'hc2903352} /* (17, 28, 21) {real, imag} */,
  {32'h42029686, 32'hc2102d8a} /* (17, 28, 20) {real, imag} */,
  {32'hc1ea213c, 32'hc007ff30} /* (17, 28, 19) {real, imag} */,
  {32'hc2289712, 32'h421e3766} /* (17, 28, 18) {real, imag} */,
  {32'h41bfa640, 32'h414cb87a} /* (17, 28, 17) {real, imag} */,
  {32'hc1aa09f0, 32'h00000000} /* (17, 28, 16) {real, imag} */,
  {32'h41bfa640, 32'hc14cb87a} /* (17, 28, 15) {real, imag} */,
  {32'hc2289712, 32'hc21e3766} /* (17, 28, 14) {real, imag} */,
  {32'hc1ea213c, 32'h4007ff30} /* (17, 28, 13) {real, imag} */,
  {32'h42029686, 32'h42102d8a} /* (17, 28, 12) {real, imag} */,
  {32'h42592726, 32'h42903352} /* (17, 28, 11) {real, imag} */,
  {32'h4185858f, 32'hc1048348} /* (17, 28, 10) {real, imag} */,
  {32'h42820c4a, 32'hc1fb97e1} /* (17, 28, 9) {real, imag} */,
  {32'h41bbcf82, 32'h41c6b734} /* (17, 28, 8) {real, imag} */,
  {32'hc0fe3508, 32'h4215e397} /* (17, 28, 7) {real, imag} */,
  {32'h430ab31d, 32'hc113387a} /* (17, 28, 6) {real, imag} */,
  {32'h430b90b6, 32'h425211ec} /* (17, 28, 5) {real, imag} */,
  {32'hc3261405, 32'hc26b8e36} /* (17, 28, 4) {real, imag} */,
  {32'hc160cd28, 32'h41a8bce7} /* (17, 28, 3) {real, imag} */,
  {32'h4482c906, 32'h43cf5d1a} /* (17, 28, 2) {real, imag} */,
  {32'hc549b455, 32'hc413a116} /* (17, 28, 1) {real, imag} */,
  {32'hc532fd44, 32'h00000000} /* (17, 28, 0) {real, imag} */,
  {32'hc5485a97, 32'h43ca91b0} /* (17, 27, 31) {real, imag} */,
  {32'h448e1bec, 32'hc3fb8640} /* (17, 27, 30) {real, imag} */,
  {32'hc29c4d4c, 32'hc2982448} /* (17, 27, 29) {real, imag} */,
  {32'hc36f6663, 32'h4355609b} /* (17, 27, 28) {real, imag} */,
  {32'h43269661, 32'hc2818300} /* (17, 27, 27) {real, imag} */,
  {32'h42a0b19d, 32'h4295784d} /* (17, 27, 26) {real, imag} */,
  {32'hc0802130, 32'hc0839060} /* (17, 27, 25) {real, imag} */,
  {32'h42e4de15, 32'hc16a37b8} /* (17, 27, 24) {real, imag} */,
  {32'h42e6efa0, 32'hc21190d9} /* (17, 27, 23) {real, imag} */,
  {32'h40878b90, 32'hc1b9ae24} /* (17, 27, 22) {real, imag} */,
  {32'h42aed4e4, 32'hc2a5d49f} /* (17, 27, 21) {real, imag} */,
  {32'h42a93fc8, 32'h42412a66} /* (17, 27, 20) {real, imag} */,
  {32'h420d7c0d, 32'h423e3b83} /* (17, 27, 19) {real, imag} */,
  {32'hc20e2494, 32'hc25cc7f8} /* (17, 27, 18) {real, imag} */,
  {32'h41b86bc4, 32'h42a2d629} /* (17, 27, 17) {real, imag} */,
  {32'h4179036c, 32'h00000000} /* (17, 27, 16) {real, imag} */,
  {32'h41b86bc4, 32'hc2a2d629} /* (17, 27, 15) {real, imag} */,
  {32'hc20e2494, 32'h425cc7f8} /* (17, 27, 14) {real, imag} */,
  {32'h420d7c0d, 32'hc23e3b83} /* (17, 27, 13) {real, imag} */,
  {32'h42a93fc8, 32'hc2412a66} /* (17, 27, 12) {real, imag} */,
  {32'h42aed4e4, 32'h42a5d49f} /* (17, 27, 11) {real, imag} */,
  {32'h40878b90, 32'h41b9ae24} /* (17, 27, 10) {real, imag} */,
  {32'h42e6efa0, 32'h421190d9} /* (17, 27, 9) {real, imag} */,
  {32'h42e4de15, 32'h416a37b8} /* (17, 27, 8) {real, imag} */,
  {32'hc0802130, 32'h40839060} /* (17, 27, 7) {real, imag} */,
  {32'h42a0b19d, 32'hc295784d} /* (17, 27, 6) {real, imag} */,
  {32'h43269661, 32'h42818300} /* (17, 27, 5) {real, imag} */,
  {32'hc36f6663, 32'hc355609b} /* (17, 27, 4) {real, imag} */,
  {32'hc29c4d4c, 32'h42982448} /* (17, 27, 3) {real, imag} */,
  {32'h448e1bec, 32'h43fb8640} /* (17, 27, 2) {real, imag} */,
  {32'hc5485a97, 32'hc3ca91b0} /* (17, 27, 1) {real, imag} */,
  {32'hc539a72c, 32'h00000000} /* (17, 27, 0) {real, imag} */,
  {32'hc536c6ed, 32'h435e930c} /* (17, 26, 31) {real, imag} */,
  {32'h44863e36, 32'hc3d983a2} /* (17, 26, 30) {real, imag} */,
  {32'hc1ff52aa, 32'h411b2fae} /* (17, 26, 29) {real, imag} */,
  {32'hc38aa62a, 32'hc2899e88} /* (17, 26, 28) {real, imag} */,
  {32'h431b4574, 32'hc2105f0a} /* (17, 26, 27) {real, imag} */,
  {32'hc147eee8, 32'h41aa3c5a} /* (17, 26, 26) {real, imag} */,
  {32'hc1e3ddc3, 32'h42847b48} /* (17, 26, 25) {real, imag} */,
  {32'h42a5a7d9, 32'hc20ae5b0} /* (17, 26, 24) {real, imag} */,
  {32'h401f6284, 32'hc2b7098c} /* (17, 26, 23) {real, imag} */,
  {32'hc18d836e, 32'h41710160} /* (17, 26, 22) {real, imag} */,
  {32'hbfaa6b40, 32'hc24d9663} /* (17, 26, 21) {real, imag} */,
  {32'h41ca36b1, 32'h429bde85} /* (17, 26, 20) {real, imag} */,
  {32'hc26983a5, 32'hc269db0c} /* (17, 26, 19) {real, imag} */,
  {32'h42078993, 32'hc23a5a38} /* (17, 26, 18) {real, imag} */,
  {32'hc0ce3840, 32'h420f6928} /* (17, 26, 17) {real, imag} */,
  {32'hc2a2ad36, 32'h00000000} /* (17, 26, 16) {real, imag} */,
  {32'hc0ce3840, 32'hc20f6928} /* (17, 26, 15) {real, imag} */,
  {32'h42078993, 32'h423a5a38} /* (17, 26, 14) {real, imag} */,
  {32'hc26983a5, 32'h4269db0c} /* (17, 26, 13) {real, imag} */,
  {32'h41ca36b1, 32'hc29bde85} /* (17, 26, 12) {real, imag} */,
  {32'hbfaa6b40, 32'h424d9663} /* (17, 26, 11) {real, imag} */,
  {32'hc18d836e, 32'hc1710160} /* (17, 26, 10) {real, imag} */,
  {32'h401f6284, 32'h42b7098c} /* (17, 26, 9) {real, imag} */,
  {32'h42a5a7d9, 32'h420ae5b0} /* (17, 26, 8) {real, imag} */,
  {32'hc1e3ddc3, 32'hc2847b48} /* (17, 26, 7) {real, imag} */,
  {32'hc147eee8, 32'hc1aa3c5a} /* (17, 26, 6) {real, imag} */,
  {32'h431b4574, 32'h42105f0a} /* (17, 26, 5) {real, imag} */,
  {32'hc38aa62a, 32'h42899e88} /* (17, 26, 4) {real, imag} */,
  {32'hc1ff52aa, 32'hc11b2fae} /* (17, 26, 3) {real, imag} */,
  {32'h44863e36, 32'h43d983a2} /* (17, 26, 2) {real, imag} */,
  {32'hc536c6ed, 32'hc35e930c} /* (17, 26, 1) {real, imag} */,
  {32'hc5341ed8, 32'h00000000} /* (17, 26, 0) {real, imag} */,
  {32'hc52d0265, 32'h433a0450} /* (17, 25, 31) {real, imag} */,
  {32'h4462a15b, 32'hc3913080} /* (17, 25, 30) {real, imag} */,
  {32'hc16a0a64, 32'hc20c734c} /* (17, 25, 29) {real, imag} */,
  {32'hc395efc8, 32'hc295e1ae} /* (17, 25, 28) {real, imag} */,
  {32'h434d33a7, 32'hc2a05907} /* (17, 25, 27) {real, imag} */,
  {32'h428d40c4, 32'hc2246e98} /* (17, 25, 26) {real, imag} */,
  {32'hc2cfbaa6, 32'h4195d318} /* (17, 25, 25) {real, imag} */,
  {32'h434c7dc4, 32'hc3191f6e} /* (17, 25, 24) {real, imag} */,
  {32'h418cdea0, 32'h422d4989} /* (17, 25, 23) {real, imag} */,
  {32'hc18c7c4a, 32'hc1c7bf23} /* (17, 25, 22) {real, imag} */,
  {32'h411e14b5, 32'hc272fd40} /* (17, 25, 21) {real, imag} */,
  {32'h40d690fe, 32'hc191aeea} /* (17, 25, 20) {real, imag} */,
  {32'hc26c3a14, 32'hc206a02a} /* (17, 25, 19) {real, imag} */,
  {32'h41d23462, 32'hc28ce112} /* (17, 25, 18) {real, imag} */,
  {32'h40a34df1, 32'h40745620} /* (17, 25, 17) {real, imag} */,
  {32'hc1ac9c20, 32'h00000000} /* (17, 25, 16) {real, imag} */,
  {32'h40a34df1, 32'hc0745620} /* (17, 25, 15) {real, imag} */,
  {32'h41d23462, 32'h428ce112} /* (17, 25, 14) {real, imag} */,
  {32'hc26c3a14, 32'h4206a02a} /* (17, 25, 13) {real, imag} */,
  {32'h40d690fe, 32'h4191aeea} /* (17, 25, 12) {real, imag} */,
  {32'h411e14b5, 32'h4272fd40} /* (17, 25, 11) {real, imag} */,
  {32'hc18c7c4a, 32'h41c7bf23} /* (17, 25, 10) {real, imag} */,
  {32'h418cdea0, 32'hc22d4989} /* (17, 25, 9) {real, imag} */,
  {32'h434c7dc4, 32'h43191f6e} /* (17, 25, 8) {real, imag} */,
  {32'hc2cfbaa6, 32'hc195d318} /* (17, 25, 7) {real, imag} */,
  {32'h428d40c4, 32'h42246e98} /* (17, 25, 6) {real, imag} */,
  {32'h434d33a7, 32'h42a05907} /* (17, 25, 5) {real, imag} */,
  {32'hc395efc8, 32'h4295e1ae} /* (17, 25, 4) {real, imag} */,
  {32'hc16a0a64, 32'h420c734c} /* (17, 25, 3) {real, imag} */,
  {32'h4462a15b, 32'h43913080} /* (17, 25, 2) {real, imag} */,
  {32'hc52d0265, 32'hc33a0450} /* (17, 25, 1) {real, imag} */,
  {32'hc5267050, 32'h00000000} /* (17, 25, 0) {real, imag} */,
  {32'hc51bd1a1, 32'h4313a3aa} /* (17, 24, 31) {real, imag} */,
  {32'h446eebca, 32'hc2d06dc8} /* (17, 24, 30) {real, imag} */,
  {32'hc2573c2b, 32'hc28c6d8b} /* (17, 24, 29) {real, imag} */,
  {32'hc3a41372, 32'hc2855d47} /* (17, 24, 28) {real, imag} */,
  {32'h438d1d00, 32'hc34e9952} /* (17, 24, 27) {real, imag} */,
  {32'hc27b5dfc, 32'hc280e818} /* (17, 24, 26) {real, imag} */,
  {32'hc2756b66, 32'h41fc43df} /* (17, 24, 25) {real, imag} */,
  {32'h438ba308, 32'h3fd34960} /* (17, 24, 24) {real, imag} */,
  {32'hc28b614b, 32'hc2514fa8} /* (17, 24, 23) {real, imag} */,
  {32'hbf6a5580, 32'h423e24ce} /* (17, 24, 22) {real, imag} */,
  {32'h4264146a, 32'hc2f0b728} /* (17, 24, 21) {real, imag} */,
  {32'hc26061e2, 32'hc0dd2930} /* (17, 24, 20) {real, imag} */,
  {32'h42650844, 32'hc20598de} /* (17, 24, 19) {real, imag} */,
  {32'h40884fe7, 32'hc2ea6ea4} /* (17, 24, 18) {real, imag} */,
  {32'h42255e6a, 32'hc092a828} /* (17, 24, 17) {real, imag} */,
  {32'hc2eb9f86, 32'h00000000} /* (17, 24, 16) {real, imag} */,
  {32'h42255e6a, 32'h4092a828} /* (17, 24, 15) {real, imag} */,
  {32'h40884fe7, 32'h42ea6ea4} /* (17, 24, 14) {real, imag} */,
  {32'h42650844, 32'h420598de} /* (17, 24, 13) {real, imag} */,
  {32'hc26061e2, 32'h40dd2930} /* (17, 24, 12) {real, imag} */,
  {32'h4264146a, 32'h42f0b728} /* (17, 24, 11) {real, imag} */,
  {32'hbf6a5580, 32'hc23e24ce} /* (17, 24, 10) {real, imag} */,
  {32'hc28b614b, 32'h42514fa8} /* (17, 24, 9) {real, imag} */,
  {32'h438ba308, 32'hbfd34960} /* (17, 24, 8) {real, imag} */,
  {32'hc2756b66, 32'hc1fc43df} /* (17, 24, 7) {real, imag} */,
  {32'hc27b5dfc, 32'h4280e818} /* (17, 24, 6) {real, imag} */,
  {32'h438d1d00, 32'h434e9952} /* (17, 24, 5) {real, imag} */,
  {32'hc3a41372, 32'h42855d47} /* (17, 24, 4) {real, imag} */,
  {32'hc2573c2b, 32'h428c6d8b} /* (17, 24, 3) {real, imag} */,
  {32'h446eebca, 32'h42d06dc8} /* (17, 24, 2) {real, imag} */,
  {32'hc51bd1a1, 32'hc313a3aa} /* (17, 24, 1) {real, imag} */,
  {32'hc52119f2, 32'h00000000} /* (17, 24, 0) {real, imag} */,
  {32'hc502a5b2, 32'h42cd63fc} /* (17, 23, 31) {real, imag} */,
  {32'h445cbc47, 32'hc29026d3} /* (17, 23, 30) {real, imag} */,
  {32'h42973eb6, 32'h416192c4} /* (17, 23, 29) {real, imag} */,
  {32'hc30a1cac, 32'hc2b4e9f6} /* (17, 23, 28) {real, imag} */,
  {32'h43628513, 32'hc3153120} /* (17, 23, 27) {real, imag} */,
  {32'hc1fc3828, 32'hc2cbc754} /* (17, 23, 26) {real, imag} */,
  {32'hc1d80864, 32'hbf850780} /* (17, 23, 25) {real, imag} */,
  {32'h428d461b, 32'hc2075e82} /* (17, 23, 24) {real, imag} */,
  {32'hc1870360, 32'hc26228f4} /* (17, 23, 23) {real, imag} */,
  {32'hc1cd920a, 32'h4287722a} /* (17, 23, 22) {real, imag} */,
  {32'hc1caf3ba, 32'h42db51f4} /* (17, 23, 21) {real, imag} */,
  {32'h4196cea6, 32'hc187cb7c} /* (17, 23, 20) {real, imag} */,
  {32'h41d1b28b, 32'h40fde608} /* (17, 23, 19) {real, imag} */,
  {32'hc24a69f8, 32'hc1903dc0} /* (17, 23, 18) {real, imag} */,
  {32'h4202a77c, 32'h4231ea48} /* (17, 23, 17) {real, imag} */,
  {32'h41bd31db, 32'h00000000} /* (17, 23, 16) {real, imag} */,
  {32'h4202a77c, 32'hc231ea48} /* (17, 23, 15) {real, imag} */,
  {32'hc24a69f8, 32'h41903dc0} /* (17, 23, 14) {real, imag} */,
  {32'h41d1b28b, 32'hc0fde608} /* (17, 23, 13) {real, imag} */,
  {32'h4196cea6, 32'h4187cb7c} /* (17, 23, 12) {real, imag} */,
  {32'hc1caf3ba, 32'hc2db51f4} /* (17, 23, 11) {real, imag} */,
  {32'hc1cd920a, 32'hc287722a} /* (17, 23, 10) {real, imag} */,
  {32'hc1870360, 32'h426228f4} /* (17, 23, 9) {real, imag} */,
  {32'h428d461b, 32'h42075e82} /* (17, 23, 8) {real, imag} */,
  {32'hc1d80864, 32'h3f850780} /* (17, 23, 7) {real, imag} */,
  {32'hc1fc3828, 32'h42cbc754} /* (17, 23, 6) {real, imag} */,
  {32'h43628513, 32'h43153120} /* (17, 23, 5) {real, imag} */,
  {32'hc30a1cac, 32'h42b4e9f6} /* (17, 23, 4) {real, imag} */,
  {32'h42973eb6, 32'hc16192c4} /* (17, 23, 3) {real, imag} */,
  {32'h445cbc47, 32'h429026d3} /* (17, 23, 2) {real, imag} */,
  {32'hc502a5b2, 32'hc2cd63fc} /* (17, 23, 1) {real, imag} */,
  {32'hc506929d, 32'h00000000} /* (17, 23, 0) {real, imag} */,
  {32'hc4b6a6f2, 32'h42fd9fc8} /* (17, 22, 31) {real, imag} */,
  {32'h44222d97, 32'hc2fdff52} /* (17, 22, 30) {real, imag} */,
  {32'hc28e5dd4, 32'hc0882e98} /* (17, 22, 29) {real, imag} */,
  {32'hc2e48000, 32'h41df477c} /* (17, 22, 28) {real, imag} */,
  {32'h42dd4116, 32'hc2f7cc4b} /* (17, 22, 27) {real, imag} */,
  {32'hc1f715fc, 32'h41645de8} /* (17, 22, 26) {real, imag} */,
  {32'hc271f071, 32'h42268e6e} /* (17, 22, 25) {real, imag} */,
  {32'h41cf14f0, 32'hc2866dc1} /* (17, 22, 24) {real, imag} */,
  {32'h422e37a6, 32'hc1641454} /* (17, 22, 23) {real, imag} */,
  {32'hc1dcb172, 32'h42717a8e} /* (17, 22, 22) {real, imag} */,
  {32'h43046cb2, 32'hbf1570c0} /* (17, 22, 21) {real, imag} */,
  {32'h417672b0, 32'h4204422c} /* (17, 22, 20) {real, imag} */,
  {32'h403e0d70, 32'hc03a41b0} /* (17, 22, 19) {real, imag} */,
  {32'hc16aec98, 32'hc205fb66} /* (17, 22, 18) {real, imag} */,
  {32'hc0e8c940, 32'h422f164b} /* (17, 22, 17) {real, imag} */,
  {32'hc26bf93b, 32'h00000000} /* (17, 22, 16) {real, imag} */,
  {32'hc0e8c940, 32'hc22f164b} /* (17, 22, 15) {real, imag} */,
  {32'hc16aec98, 32'h4205fb66} /* (17, 22, 14) {real, imag} */,
  {32'h403e0d70, 32'h403a41b0} /* (17, 22, 13) {real, imag} */,
  {32'h417672b0, 32'hc204422c} /* (17, 22, 12) {real, imag} */,
  {32'h43046cb2, 32'h3f1570c0} /* (17, 22, 11) {real, imag} */,
  {32'hc1dcb172, 32'hc2717a8e} /* (17, 22, 10) {real, imag} */,
  {32'h422e37a6, 32'h41641454} /* (17, 22, 9) {real, imag} */,
  {32'h41cf14f0, 32'h42866dc1} /* (17, 22, 8) {real, imag} */,
  {32'hc271f071, 32'hc2268e6e} /* (17, 22, 7) {real, imag} */,
  {32'hc1f715fc, 32'hc1645de8} /* (17, 22, 6) {real, imag} */,
  {32'h42dd4116, 32'h42f7cc4b} /* (17, 22, 5) {real, imag} */,
  {32'hc2e48000, 32'hc1df477c} /* (17, 22, 4) {real, imag} */,
  {32'hc28e5dd4, 32'h40882e98} /* (17, 22, 3) {real, imag} */,
  {32'h44222d97, 32'h42fdff52} /* (17, 22, 2) {real, imag} */,
  {32'hc4b6a6f2, 32'hc2fd9fc8} /* (17, 22, 1) {real, imag} */,
  {32'hc4c53cf2, 32'h00000000} /* (17, 22, 0) {real, imag} */,
  {32'hc413be73, 32'h43423bf8} /* (17, 21, 31) {real, imag} */,
  {32'h437ee008, 32'h4320e656} /* (17, 21, 30) {real, imag} */,
  {32'hc211387c, 32'h42037dd8} /* (17, 21, 29) {real, imag} */,
  {32'hc1b9e563, 32'hc1256bd8} /* (17, 21, 28) {real, imag} */,
  {32'h42aa7e9f, 32'hc29738f3} /* (17, 21, 27) {real, imag} */,
  {32'hc1b9ae31, 32'hc22b94da} /* (17, 21, 26) {real, imag} */,
  {32'h404213c0, 32'h42e3b12f} /* (17, 21, 25) {real, imag} */,
  {32'h422bab7d, 32'hc11c9d20} /* (17, 21, 24) {real, imag} */,
  {32'h421f4e9c, 32'h4016109a} /* (17, 21, 23) {real, imag} */,
  {32'hc136d078, 32'hc2863d3a} /* (17, 21, 22) {real, imag} */,
  {32'hc193b302, 32'hc2fc4d5a} /* (17, 21, 21) {real, imag} */,
  {32'hc2200c06, 32'hc206c857} /* (17, 21, 20) {real, imag} */,
  {32'h41dce098, 32'h4030901e} /* (17, 21, 19) {real, imag} */,
  {32'hbffaeb00, 32'hbfb715e0} /* (17, 21, 18) {real, imag} */,
  {32'hc1336ecb, 32'h41979fd5} /* (17, 21, 17) {real, imag} */,
  {32'hc26c9c49, 32'h00000000} /* (17, 21, 16) {real, imag} */,
  {32'hc1336ecb, 32'hc1979fd5} /* (17, 21, 15) {real, imag} */,
  {32'hbffaeb00, 32'h3fb715e0} /* (17, 21, 14) {real, imag} */,
  {32'h41dce098, 32'hc030901e} /* (17, 21, 13) {real, imag} */,
  {32'hc2200c06, 32'h4206c857} /* (17, 21, 12) {real, imag} */,
  {32'hc193b302, 32'h42fc4d5a} /* (17, 21, 11) {real, imag} */,
  {32'hc136d078, 32'h42863d3a} /* (17, 21, 10) {real, imag} */,
  {32'h421f4e9c, 32'hc016109a} /* (17, 21, 9) {real, imag} */,
  {32'h422bab7d, 32'h411c9d20} /* (17, 21, 8) {real, imag} */,
  {32'h404213c0, 32'hc2e3b12f} /* (17, 21, 7) {real, imag} */,
  {32'hc1b9ae31, 32'h422b94da} /* (17, 21, 6) {real, imag} */,
  {32'h42aa7e9f, 32'h429738f3} /* (17, 21, 5) {real, imag} */,
  {32'hc1b9e563, 32'h41256bd8} /* (17, 21, 4) {real, imag} */,
  {32'hc211387c, 32'hc2037dd8} /* (17, 21, 3) {real, imag} */,
  {32'h437ee008, 32'hc320e656} /* (17, 21, 2) {real, imag} */,
  {32'hc413be73, 32'hc3423bf8} /* (17, 21, 1) {real, imag} */,
  {32'hc4493ea5, 32'h00000000} /* (17, 21, 0) {real, imag} */,
  {32'h44082723, 32'h429a8d24} /* (17, 20, 31) {real, imag} */,
  {32'hc38e11b5, 32'h43951656} /* (17, 20, 30) {real, imag} */,
  {32'h420eaeb0, 32'hc2e2e051} /* (17, 20, 29) {real, imag} */,
  {32'h433d9a18, 32'hc2599f0c} /* (17, 20, 28) {real, imag} */,
  {32'hc23a6faa, 32'hc26a2e6c} /* (17, 20, 27) {real, imag} */,
  {32'h41a3cabc, 32'hc2494b87} /* (17, 20, 26) {real, imag} */,
  {32'h4268d301, 32'h422271d4} /* (17, 20, 25) {real, imag} */,
  {32'hc2c63bb6, 32'h41d6de60} /* (17, 20, 24) {real, imag} */,
  {32'hc225a188, 32'hc089c304} /* (17, 20, 23) {real, imag} */,
  {32'hc24364d0, 32'hc2e8d26c} /* (17, 20, 22) {real, imag} */,
  {32'hc28dcdb0, 32'h42c288a1} /* (17, 20, 21) {real, imag} */,
  {32'h41628222, 32'h42759382} /* (17, 20, 20) {real, imag} */,
  {32'hc0d5c062, 32'h41099d14} /* (17, 20, 19) {real, imag} */,
  {32'hc2631dac, 32'h42a12ffb} /* (17, 20, 18) {real, imag} */,
  {32'h4288eff9, 32'h41f2a65b} /* (17, 20, 17) {real, imag} */,
  {32'hc0c571a1, 32'h00000000} /* (17, 20, 16) {real, imag} */,
  {32'h4288eff9, 32'hc1f2a65b} /* (17, 20, 15) {real, imag} */,
  {32'hc2631dac, 32'hc2a12ffb} /* (17, 20, 14) {real, imag} */,
  {32'hc0d5c062, 32'hc1099d14} /* (17, 20, 13) {real, imag} */,
  {32'h41628222, 32'hc2759382} /* (17, 20, 12) {real, imag} */,
  {32'hc28dcdb0, 32'hc2c288a1} /* (17, 20, 11) {real, imag} */,
  {32'hc24364d0, 32'h42e8d26c} /* (17, 20, 10) {real, imag} */,
  {32'hc225a188, 32'h4089c304} /* (17, 20, 9) {real, imag} */,
  {32'hc2c63bb6, 32'hc1d6de60} /* (17, 20, 8) {real, imag} */,
  {32'h4268d301, 32'hc22271d4} /* (17, 20, 7) {real, imag} */,
  {32'h41a3cabc, 32'h42494b87} /* (17, 20, 6) {real, imag} */,
  {32'hc23a6faa, 32'h426a2e6c} /* (17, 20, 5) {real, imag} */,
  {32'h433d9a18, 32'h42599f0c} /* (17, 20, 4) {real, imag} */,
  {32'h420eaeb0, 32'h42e2e051} /* (17, 20, 3) {real, imag} */,
  {32'hc38e11b5, 32'hc3951656} /* (17, 20, 2) {real, imag} */,
  {32'h44082723, 32'hc29a8d24} /* (17, 20, 1) {real, imag} */,
  {32'h434a9a04, 32'h00000000} /* (17, 20, 0) {real, imag} */,
  {32'h44b0507e, 32'hc32b9e52} /* (17, 19, 31) {real, imag} */,
  {32'hc412c24a, 32'h439bbd16} /* (17, 19, 30) {real, imag} */,
  {32'h4301c857, 32'h42cdbe76} /* (17, 19, 29) {real, imag} */,
  {32'h435c6bb2, 32'hc1e21baa} /* (17, 19, 28) {real, imag} */,
  {32'hc2d59792, 32'h41e512c4} /* (17, 19, 27) {real, imag} */,
  {32'hc2b7d8c2, 32'h421eeff4} /* (17, 19, 26) {real, imag} */,
  {32'h425d7a48, 32'hc27feb64} /* (17, 19, 25) {real, imag} */,
  {32'h42321950, 32'h42fb6416} /* (17, 19, 24) {real, imag} */,
  {32'hc240598a, 32'h420af076} /* (17, 19, 23) {real, imag} */,
  {32'h40e661d8, 32'h42ada6cf} /* (17, 19, 22) {real, imag} */,
  {32'h41c70dec, 32'h416b2bdc} /* (17, 19, 21) {real, imag} */,
  {32'h422a9ffc, 32'h400bdda0} /* (17, 19, 20) {real, imag} */,
  {32'h42055047, 32'h4227926a} /* (17, 19, 19) {real, imag} */,
  {32'h4210bb41, 32'hc198994c} /* (17, 19, 18) {real, imag} */,
  {32'h40c992c0, 32'hc2509132} /* (17, 19, 17) {real, imag} */,
  {32'hc2492a1c, 32'h00000000} /* (17, 19, 16) {real, imag} */,
  {32'h40c992c0, 32'h42509132} /* (17, 19, 15) {real, imag} */,
  {32'h4210bb41, 32'h4198994c} /* (17, 19, 14) {real, imag} */,
  {32'h42055047, 32'hc227926a} /* (17, 19, 13) {real, imag} */,
  {32'h422a9ffc, 32'hc00bdda0} /* (17, 19, 12) {real, imag} */,
  {32'h41c70dec, 32'hc16b2bdc} /* (17, 19, 11) {real, imag} */,
  {32'h40e661d8, 32'hc2ada6cf} /* (17, 19, 10) {real, imag} */,
  {32'hc240598a, 32'hc20af076} /* (17, 19, 9) {real, imag} */,
  {32'h42321950, 32'hc2fb6416} /* (17, 19, 8) {real, imag} */,
  {32'h425d7a48, 32'h427feb64} /* (17, 19, 7) {real, imag} */,
  {32'hc2b7d8c2, 32'hc21eeff4} /* (17, 19, 6) {real, imag} */,
  {32'hc2d59792, 32'hc1e512c4} /* (17, 19, 5) {real, imag} */,
  {32'h435c6bb2, 32'h41e21baa} /* (17, 19, 4) {real, imag} */,
  {32'h4301c857, 32'hc2cdbe76} /* (17, 19, 3) {real, imag} */,
  {32'hc412c24a, 32'hc39bbd16} /* (17, 19, 2) {real, imag} */,
  {32'h44b0507e, 32'h432b9e52} /* (17, 19, 1) {real, imag} */,
  {32'h44558985, 32'h00000000} /* (17, 19, 0) {real, imag} */,
  {32'h44f6ea8b, 32'hc2985a5c} /* (17, 18, 31) {real, imag} */,
  {32'hc446fae7, 32'h43103e86} /* (17, 18, 30) {real, imag} */,
  {32'h431b9db6, 32'h42607688} /* (17, 18, 29) {real, imag} */,
  {32'h4383997b, 32'hc125c120} /* (17, 18, 28) {real, imag} */,
  {32'hc3882440, 32'h43373e44} /* (17, 18, 27) {real, imag} */,
  {32'hc30a09ab, 32'h42449394} /* (17, 18, 26) {real, imag} */,
  {32'h42b1a52d, 32'hc1bfffe9} /* (17, 18, 25) {real, imag} */,
  {32'h41bd5a7e, 32'h43414130} /* (17, 18, 24) {real, imag} */,
  {32'hc2939512, 32'hc1db2648} /* (17, 18, 23) {real, imag} */,
  {32'h424d27f3, 32'hc25248e4} /* (17, 18, 22) {real, imag} */,
  {32'h4280a3b7, 32'h42885f24} /* (17, 18, 21) {real, imag} */,
  {32'hc2a9799e, 32'hc1d71ed3} /* (17, 18, 20) {real, imag} */,
  {32'h4159e09f, 32'hc21fe472} /* (17, 18, 19) {real, imag} */,
  {32'h4223c847, 32'hc23403ce} /* (17, 18, 18) {real, imag} */,
  {32'hc276f822, 32'hc2b037a3} /* (17, 18, 17) {real, imag} */,
  {32'h428409b7, 32'h00000000} /* (17, 18, 16) {real, imag} */,
  {32'hc276f822, 32'h42b037a3} /* (17, 18, 15) {real, imag} */,
  {32'h4223c847, 32'h423403ce} /* (17, 18, 14) {real, imag} */,
  {32'h4159e09f, 32'h421fe472} /* (17, 18, 13) {real, imag} */,
  {32'hc2a9799e, 32'h41d71ed3} /* (17, 18, 12) {real, imag} */,
  {32'h4280a3b7, 32'hc2885f24} /* (17, 18, 11) {real, imag} */,
  {32'h424d27f3, 32'h425248e4} /* (17, 18, 10) {real, imag} */,
  {32'hc2939512, 32'h41db2648} /* (17, 18, 9) {real, imag} */,
  {32'h41bd5a7e, 32'hc3414130} /* (17, 18, 8) {real, imag} */,
  {32'h42b1a52d, 32'h41bfffe9} /* (17, 18, 7) {real, imag} */,
  {32'hc30a09ab, 32'hc2449394} /* (17, 18, 6) {real, imag} */,
  {32'hc3882440, 32'hc3373e44} /* (17, 18, 5) {real, imag} */,
  {32'h4383997b, 32'h4125c120} /* (17, 18, 4) {real, imag} */,
  {32'h431b9db6, 32'hc2607688} /* (17, 18, 3) {real, imag} */,
  {32'hc446fae7, 32'hc3103e86} /* (17, 18, 2) {real, imag} */,
  {32'h44f6ea8b, 32'h42985a5c} /* (17, 18, 1) {real, imag} */,
  {32'h44b89718, 32'h00000000} /* (17, 18, 0) {real, imag} */,
  {32'h4509c7bf, 32'hc26f1a88} /* (17, 17, 31) {real, imag} */,
  {32'hc4881b14, 32'h42855c48} /* (17, 17, 30) {real, imag} */,
  {32'h4370843e, 32'hc2788e00} /* (17, 17, 29) {real, imag} */,
  {32'h43865f67, 32'hc1a2b3c4} /* (17, 17, 28) {real, imag} */,
  {32'hc3980553, 32'h43010dd2} /* (17, 17, 27) {real, imag} */,
  {32'hc30721ff, 32'hc2a53c66} /* (17, 17, 26) {real, imag} */,
  {32'h42c7fa53, 32'h41b87623} /* (17, 17, 25) {real, imag} */,
  {32'hc23d3c50, 32'h424bfcc6} /* (17, 17, 24) {real, imag} */,
  {32'hc0bdda28, 32'h40cb19a4} /* (17, 17, 23) {real, imag} */,
  {32'hc1dbc2b4, 32'h42841422} /* (17, 17, 22) {real, imag} */,
  {32'hc23a1e73, 32'h41d9ab04} /* (17, 17, 21) {real, imag} */,
  {32'hc097ae94, 32'hc3009b53} /* (17, 17, 20) {real, imag} */,
  {32'h42d7c057, 32'h42085f2d} /* (17, 17, 19) {real, imag} */,
  {32'hc232dad2, 32'h429d594d} /* (17, 17, 18) {real, imag} */,
  {32'h41312ccc, 32'hbfe42720} /* (17, 17, 17) {real, imag} */,
  {32'h42698b5a, 32'h00000000} /* (17, 17, 16) {real, imag} */,
  {32'h41312ccc, 32'h3fe42720} /* (17, 17, 15) {real, imag} */,
  {32'hc232dad2, 32'hc29d594d} /* (17, 17, 14) {real, imag} */,
  {32'h42d7c057, 32'hc2085f2d} /* (17, 17, 13) {real, imag} */,
  {32'hc097ae94, 32'h43009b53} /* (17, 17, 12) {real, imag} */,
  {32'hc23a1e73, 32'hc1d9ab04} /* (17, 17, 11) {real, imag} */,
  {32'hc1dbc2b4, 32'hc2841422} /* (17, 17, 10) {real, imag} */,
  {32'hc0bdda28, 32'hc0cb19a4} /* (17, 17, 9) {real, imag} */,
  {32'hc23d3c50, 32'hc24bfcc6} /* (17, 17, 8) {real, imag} */,
  {32'h42c7fa53, 32'hc1b87623} /* (17, 17, 7) {real, imag} */,
  {32'hc30721ff, 32'h42a53c66} /* (17, 17, 6) {real, imag} */,
  {32'hc3980553, 32'hc3010dd2} /* (17, 17, 5) {real, imag} */,
  {32'h43865f67, 32'h41a2b3c4} /* (17, 17, 4) {real, imag} */,
  {32'h4370843e, 32'h42788e00} /* (17, 17, 3) {real, imag} */,
  {32'hc4881b14, 32'hc2855c48} /* (17, 17, 2) {real, imag} */,
  {32'h4509c7bf, 32'h426f1a88} /* (17, 17, 1) {real, imag} */,
  {32'h44e193d6, 32'h00000000} /* (17, 17, 0) {real, imag} */,
  {32'h4514a63e, 32'hc323f8b0} /* (17, 16, 31) {real, imag} */,
  {32'hc49100b0, 32'h431814f8} /* (17, 16, 30) {real, imag} */,
  {32'h43200772, 32'hc31f8f7a} /* (17, 16, 29) {real, imag} */,
  {32'h4396f416, 32'h413cea8c} /* (17, 16, 28) {real, imag} */,
  {32'hc39b584b, 32'h4332e98c} /* (17, 16, 27) {real, imag} */,
  {32'h41f7555b, 32'hc292685e} /* (17, 16, 26) {real, imag} */,
  {32'h425e3a04, 32'h42324f18} /* (17, 16, 25) {real, imag} */,
  {32'hc1fdb244, 32'h426ebd45} /* (17, 16, 24) {real, imag} */,
  {32'h427460bf, 32'h40822da8} /* (17, 16, 23) {real, imag} */,
  {32'hc24fd83a, 32'h4287f6fd} /* (17, 16, 22) {real, imag} */,
  {32'h42b065b6, 32'hc174366b} /* (17, 16, 21) {real, imag} */,
  {32'hc2453334, 32'h420c7298} /* (17, 16, 20) {real, imag} */,
  {32'hc1844f79, 32'hc0c5c296} /* (17, 16, 19) {real, imag} */,
  {32'h42ba90ed, 32'h41807334} /* (17, 16, 18) {real, imag} */,
  {32'hc2d37982, 32'h42110d62} /* (17, 16, 17) {real, imag} */,
  {32'h4259a181, 32'h00000000} /* (17, 16, 16) {real, imag} */,
  {32'hc2d37982, 32'hc2110d62} /* (17, 16, 15) {real, imag} */,
  {32'h42ba90ed, 32'hc1807334} /* (17, 16, 14) {real, imag} */,
  {32'hc1844f79, 32'h40c5c296} /* (17, 16, 13) {real, imag} */,
  {32'hc2453334, 32'hc20c7298} /* (17, 16, 12) {real, imag} */,
  {32'h42b065b6, 32'h4174366b} /* (17, 16, 11) {real, imag} */,
  {32'hc24fd83a, 32'hc287f6fd} /* (17, 16, 10) {real, imag} */,
  {32'h427460bf, 32'hc0822da8} /* (17, 16, 9) {real, imag} */,
  {32'hc1fdb244, 32'hc26ebd45} /* (17, 16, 8) {real, imag} */,
  {32'h425e3a04, 32'hc2324f18} /* (17, 16, 7) {real, imag} */,
  {32'h41f7555b, 32'h4292685e} /* (17, 16, 6) {real, imag} */,
  {32'hc39b584b, 32'hc332e98c} /* (17, 16, 5) {real, imag} */,
  {32'h4396f416, 32'hc13cea8c} /* (17, 16, 4) {real, imag} */,
  {32'h43200772, 32'h431f8f7a} /* (17, 16, 3) {real, imag} */,
  {32'hc49100b0, 32'hc31814f8} /* (17, 16, 2) {real, imag} */,
  {32'h4514a63e, 32'h4323f8b0} /* (17, 16, 1) {real, imag} */,
  {32'h44cb3a74, 32'h00000000} /* (17, 16, 0) {real, imag} */,
  {32'h450ea75f, 32'hc187e170} /* (17, 15, 31) {real, imag} */,
  {32'hc486ffc0, 32'h4362f834} /* (17, 15, 30) {real, imag} */,
  {32'h42f88c69, 32'hc2d297d8} /* (17, 15, 29) {real, imag} */,
  {32'h4348271a, 32'h42749e92} /* (17, 15, 28) {real, imag} */,
  {32'hc3a66c2f, 32'h43851564} /* (17, 15, 27) {real, imag} */,
  {32'hc235874c, 32'hc35e4ed9} /* (17, 15, 26) {real, imag} */,
  {32'h42cb0b65, 32'hc0cefb9c} /* (17, 15, 25) {real, imag} */,
  {32'hc31d26be, 32'h42ad16cb} /* (17, 15, 24) {real, imag} */,
  {32'hc2a3a69a, 32'hc21b1902} /* (17, 15, 23) {real, imag} */,
  {32'h4292d136, 32'hc01fbb30} /* (17, 15, 22) {real, imag} */,
  {32'h41b3ed22, 32'h42cc079f} /* (17, 15, 21) {real, imag} */,
  {32'h4287f0d5, 32'hc20e0343} /* (17, 15, 20) {real, imag} */,
  {32'h413d7f78, 32'hc214405f} /* (17, 15, 19) {real, imag} */,
  {32'h418e7a8b, 32'h41be4121} /* (17, 15, 18) {real, imag} */,
  {32'hc02eca72, 32'hc2b31a04} /* (17, 15, 17) {real, imag} */,
  {32'h41e6000b, 32'h00000000} /* (17, 15, 16) {real, imag} */,
  {32'hc02eca72, 32'h42b31a04} /* (17, 15, 15) {real, imag} */,
  {32'h418e7a8b, 32'hc1be4121} /* (17, 15, 14) {real, imag} */,
  {32'h413d7f78, 32'h4214405f} /* (17, 15, 13) {real, imag} */,
  {32'h4287f0d5, 32'h420e0343} /* (17, 15, 12) {real, imag} */,
  {32'h41b3ed22, 32'hc2cc079f} /* (17, 15, 11) {real, imag} */,
  {32'h4292d136, 32'h401fbb30} /* (17, 15, 10) {real, imag} */,
  {32'hc2a3a69a, 32'h421b1902} /* (17, 15, 9) {real, imag} */,
  {32'hc31d26be, 32'hc2ad16cb} /* (17, 15, 8) {real, imag} */,
  {32'h42cb0b65, 32'h40cefb9c} /* (17, 15, 7) {real, imag} */,
  {32'hc235874c, 32'h435e4ed9} /* (17, 15, 6) {real, imag} */,
  {32'hc3a66c2f, 32'hc3851564} /* (17, 15, 5) {real, imag} */,
  {32'h4348271a, 32'hc2749e92} /* (17, 15, 4) {real, imag} */,
  {32'h42f88c69, 32'h42d297d8} /* (17, 15, 3) {real, imag} */,
  {32'hc486ffc0, 32'hc362f834} /* (17, 15, 2) {real, imag} */,
  {32'h450ea75f, 32'h4187e170} /* (17, 15, 1) {real, imag} */,
  {32'h44dc9a3e, 32'h00000000} /* (17, 15, 0) {real, imag} */,
  {32'h45060e09, 32'h41675e60} /* (17, 14, 31) {real, imag} */,
  {32'hc46b83c1, 32'h430ace8a} /* (17, 14, 30) {real, imag} */,
  {32'h430e95c6, 32'hc20ac680} /* (17, 14, 29) {real, imag} */,
  {32'h42d08e54, 32'h427feb28} /* (17, 14, 28) {real, imag} */,
  {32'hc3d188da, 32'h436180f6} /* (17, 14, 27) {real, imag} */,
  {32'h428b9022, 32'h428ee846} /* (17, 14, 26) {real, imag} */,
  {32'hc2a3a4bf, 32'hc203e594} /* (17, 14, 25) {real, imag} */,
  {32'hc2453995, 32'h42d3e9e1} /* (17, 14, 24) {real, imag} */,
  {32'h42944fde, 32'hc23e8674} /* (17, 14, 23) {real, imag} */,
  {32'h4242bd95, 32'h4276de14} /* (17, 14, 22) {real, imag} */,
  {32'h419ac0ab, 32'h422d0158} /* (17, 14, 21) {real, imag} */,
  {32'hc2657df4, 32'hc21fc802} /* (17, 14, 20) {real, imag} */,
  {32'h41c3be10, 32'h40dd90a8} /* (17, 14, 19) {real, imag} */,
  {32'hc217c259, 32'hc30aafae} /* (17, 14, 18) {real, imag} */,
  {32'h413102e8, 32'h419367fc} /* (17, 14, 17) {real, imag} */,
  {32'hc24cfe06, 32'h00000000} /* (17, 14, 16) {real, imag} */,
  {32'h413102e8, 32'hc19367fc} /* (17, 14, 15) {real, imag} */,
  {32'hc217c259, 32'h430aafae} /* (17, 14, 14) {real, imag} */,
  {32'h41c3be10, 32'hc0dd90a8} /* (17, 14, 13) {real, imag} */,
  {32'hc2657df4, 32'h421fc802} /* (17, 14, 12) {real, imag} */,
  {32'h419ac0ab, 32'hc22d0158} /* (17, 14, 11) {real, imag} */,
  {32'h4242bd95, 32'hc276de14} /* (17, 14, 10) {real, imag} */,
  {32'h42944fde, 32'h423e8674} /* (17, 14, 9) {real, imag} */,
  {32'hc2453995, 32'hc2d3e9e1} /* (17, 14, 8) {real, imag} */,
  {32'hc2a3a4bf, 32'h4203e594} /* (17, 14, 7) {real, imag} */,
  {32'h428b9022, 32'hc28ee846} /* (17, 14, 6) {real, imag} */,
  {32'hc3d188da, 32'hc36180f6} /* (17, 14, 5) {real, imag} */,
  {32'h42d08e54, 32'hc27feb28} /* (17, 14, 4) {real, imag} */,
  {32'h430e95c6, 32'h420ac680} /* (17, 14, 3) {real, imag} */,
  {32'hc46b83c1, 32'hc30ace8a} /* (17, 14, 2) {real, imag} */,
  {32'h45060e09, 32'hc1675e60} /* (17, 14, 1) {real, imag} */,
  {32'h44cd56ea, 32'h00000000} /* (17, 14, 0) {real, imag} */,
  {32'h44dc9050, 32'h432805d2} /* (17, 13, 31) {real, imag} */,
  {32'hc46a938e, 32'h433a1395} /* (17, 13, 30) {real, imag} */,
  {32'h4366a8e5, 32'hc2f555e6} /* (17, 13, 29) {real, imag} */,
  {32'h42263f90, 32'h4279aed7} /* (17, 13, 28) {real, imag} */,
  {32'hc36e105b, 32'h43559fac} /* (17, 13, 27) {real, imag} */,
  {32'hc0f177d8, 32'hc0339758} /* (17, 13, 26) {real, imag} */,
  {32'hc2be5054, 32'hc2514b58} /* (17, 13, 25) {real, imag} */,
  {32'h427a6e74, 32'h42bb07aa} /* (17, 13, 24) {real, imag} */,
  {32'h424a9b1c, 32'h41dfc264} /* (17, 13, 23) {real, imag} */,
  {32'h421eeae3, 32'hc1f69f17} /* (17, 13, 22) {real, imag} */,
  {32'hbff56b40, 32'hc25a279b} /* (17, 13, 21) {real, imag} */,
  {32'hc20a5788, 32'hc22aad40} /* (17, 13, 20) {real, imag} */,
  {32'h423c3cff, 32'h410fc7f2} /* (17, 13, 19) {real, imag} */,
  {32'hc12f3864, 32'hc22bc2b6} /* (17, 13, 18) {real, imag} */,
  {32'h412fd1dc, 32'hc09302b0} /* (17, 13, 17) {real, imag} */,
  {32'h42f5c082, 32'h00000000} /* (17, 13, 16) {real, imag} */,
  {32'h412fd1dc, 32'h409302b0} /* (17, 13, 15) {real, imag} */,
  {32'hc12f3864, 32'h422bc2b6} /* (17, 13, 14) {real, imag} */,
  {32'h423c3cff, 32'hc10fc7f2} /* (17, 13, 13) {real, imag} */,
  {32'hc20a5788, 32'h422aad40} /* (17, 13, 12) {real, imag} */,
  {32'hbff56b40, 32'h425a279b} /* (17, 13, 11) {real, imag} */,
  {32'h421eeae3, 32'h41f69f17} /* (17, 13, 10) {real, imag} */,
  {32'h424a9b1c, 32'hc1dfc264} /* (17, 13, 9) {real, imag} */,
  {32'h427a6e74, 32'hc2bb07aa} /* (17, 13, 8) {real, imag} */,
  {32'hc2be5054, 32'h42514b58} /* (17, 13, 7) {real, imag} */,
  {32'hc0f177d8, 32'h40339758} /* (17, 13, 6) {real, imag} */,
  {32'hc36e105b, 32'hc3559fac} /* (17, 13, 5) {real, imag} */,
  {32'h42263f90, 32'hc279aed7} /* (17, 13, 4) {real, imag} */,
  {32'h4366a8e5, 32'h42f555e6} /* (17, 13, 3) {real, imag} */,
  {32'hc46a938e, 32'hc33a1395} /* (17, 13, 2) {real, imag} */,
  {32'h44dc9050, 32'hc32805d2} /* (17, 13, 1) {real, imag} */,
  {32'h44cdb3b6, 32'h00000000} /* (17, 13, 0) {real, imag} */,
  {32'h44b52806, 32'h43268d5e} /* (17, 12, 31) {real, imag} */,
  {32'hc44b3daa, 32'h43325f06} /* (17, 12, 30) {real, imag} */,
  {32'h4378ed10, 32'h41b090cc} /* (17, 12, 29) {real, imag} */,
  {32'h4300ff42, 32'h414da128} /* (17, 12, 28) {real, imag} */,
  {32'hc32b0bfa, 32'h41eb0897} /* (17, 12, 27) {real, imag} */,
  {32'hc2c3ff6b, 32'h424a60ed} /* (17, 12, 26) {real, imag} */,
  {32'hc2587063, 32'hc326cead} /* (17, 12, 25) {real, imag} */,
  {32'hc303dffc, 32'h430317d0} /* (17, 12, 24) {real, imag} */,
  {32'h42aaef27, 32'hc230bca4} /* (17, 12, 23) {real, imag} */,
  {32'h4178434a, 32'hc2049a34} /* (17, 12, 22) {real, imag} */,
  {32'hc228556e, 32'h3f4f6f80} /* (17, 12, 21) {real, imag} */,
  {32'hc0a63054, 32'h409bb10c} /* (17, 12, 20) {real, imag} */,
  {32'h4200c4ac, 32'h41a86432} /* (17, 12, 19) {real, imag} */,
  {32'hc2812509, 32'hc1f98d34} /* (17, 12, 18) {real, imag} */,
  {32'hc2546872, 32'h427a6946} /* (17, 12, 17) {real, imag} */,
  {32'h4106ebbe, 32'h00000000} /* (17, 12, 16) {real, imag} */,
  {32'hc2546872, 32'hc27a6946} /* (17, 12, 15) {real, imag} */,
  {32'hc2812509, 32'h41f98d34} /* (17, 12, 14) {real, imag} */,
  {32'h4200c4ac, 32'hc1a86432} /* (17, 12, 13) {real, imag} */,
  {32'hc0a63054, 32'hc09bb10c} /* (17, 12, 12) {real, imag} */,
  {32'hc228556e, 32'hbf4f6f80} /* (17, 12, 11) {real, imag} */,
  {32'h4178434a, 32'h42049a34} /* (17, 12, 10) {real, imag} */,
  {32'h42aaef27, 32'h4230bca4} /* (17, 12, 9) {real, imag} */,
  {32'hc303dffc, 32'hc30317d0} /* (17, 12, 8) {real, imag} */,
  {32'hc2587063, 32'h4326cead} /* (17, 12, 7) {real, imag} */,
  {32'hc2c3ff6b, 32'hc24a60ed} /* (17, 12, 6) {real, imag} */,
  {32'hc32b0bfa, 32'hc1eb0897} /* (17, 12, 5) {real, imag} */,
  {32'h4300ff42, 32'hc14da128} /* (17, 12, 4) {real, imag} */,
  {32'h4378ed10, 32'hc1b090cc} /* (17, 12, 3) {real, imag} */,
  {32'hc44b3daa, 32'hc3325f06} /* (17, 12, 2) {real, imag} */,
  {32'h44b52806, 32'hc3268d5e} /* (17, 12, 1) {real, imag} */,
  {32'h44b1be64, 32'h00000000} /* (17, 12, 0) {real, imag} */,
  {32'h4445eac7, 32'h43a46d74} /* (17, 11, 31) {real, imag} */,
  {32'hc3e30656, 32'h434a42c8} /* (17, 11, 30) {real, imag} */,
  {32'h4331d2ff, 32'h4197c451} /* (17, 11, 29) {real, imag} */,
  {32'h4212e20e, 32'hc2a29a8e} /* (17, 11, 28) {real, imag} */,
  {32'hc2930801, 32'h42e7cc2b} /* (17, 11, 27) {real, imag} */,
  {32'hc23e3e2c, 32'hc187db8a} /* (17, 11, 26) {real, imag} */,
  {32'h42644ed3, 32'h410e8db0} /* (17, 11, 25) {real, imag} */,
  {32'hc29f4054, 32'h438d8e11} /* (17, 11, 24) {real, imag} */,
  {32'h42478408, 32'h417223ec} /* (17, 11, 23) {real, imag} */,
  {32'hc2998ab6, 32'h428a5b3e} /* (17, 11, 22) {real, imag} */,
  {32'h4264037b, 32'hc286188a} /* (17, 11, 21) {real, imag} */,
  {32'hc17f7578, 32'h417012d9} /* (17, 11, 20) {real, imag} */,
  {32'h40f6ce30, 32'h414ceae8} /* (17, 11, 19) {real, imag} */,
  {32'h428f4514, 32'h425267b4} /* (17, 11, 18) {real, imag} */,
  {32'hc1e3cf1c, 32'hc1c265fd} /* (17, 11, 17) {real, imag} */,
  {32'hc32d088b, 32'h00000000} /* (17, 11, 16) {real, imag} */,
  {32'hc1e3cf1c, 32'h41c265fd} /* (17, 11, 15) {real, imag} */,
  {32'h428f4514, 32'hc25267b4} /* (17, 11, 14) {real, imag} */,
  {32'h40f6ce30, 32'hc14ceae8} /* (17, 11, 13) {real, imag} */,
  {32'hc17f7578, 32'hc17012d9} /* (17, 11, 12) {real, imag} */,
  {32'h4264037b, 32'h4286188a} /* (17, 11, 11) {real, imag} */,
  {32'hc2998ab6, 32'hc28a5b3e} /* (17, 11, 10) {real, imag} */,
  {32'h42478408, 32'hc17223ec} /* (17, 11, 9) {real, imag} */,
  {32'hc29f4054, 32'hc38d8e11} /* (17, 11, 8) {real, imag} */,
  {32'h42644ed3, 32'hc10e8db0} /* (17, 11, 7) {real, imag} */,
  {32'hc23e3e2c, 32'h4187db8a} /* (17, 11, 6) {real, imag} */,
  {32'hc2930801, 32'hc2e7cc2b} /* (17, 11, 5) {real, imag} */,
  {32'h4212e20e, 32'h42a29a8e} /* (17, 11, 4) {real, imag} */,
  {32'h4331d2ff, 32'hc197c451} /* (17, 11, 3) {real, imag} */,
  {32'hc3e30656, 32'hc34a42c8} /* (17, 11, 2) {real, imag} */,
  {32'h4445eac7, 32'hc3a46d74} /* (17, 11, 1) {real, imag} */,
  {32'h44498ff5, 32'h00000000} /* (17, 11, 0) {real, imag} */,
  {32'hc42abf33, 32'h4404f355} /* (17, 10, 31) {real, imag} */,
  {32'h42a17488, 32'hc2281cdd} /* (17, 10, 30) {real, imag} */,
  {32'h42a5acdc, 32'h42f3c40e} /* (17, 10, 29) {real, imag} */,
  {32'hc2c86064, 32'hc2ac9e55} /* (17, 10, 28) {real, imag} */,
  {32'h420b9c1c, 32'hc08e2390} /* (17, 10, 27) {real, imag} */,
  {32'h42576b46, 32'hc095d880} /* (17, 10, 26) {real, imag} */,
  {32'h42097e23, 32'h40925464} /* (17, 10, 25) {real, imag} */,
  {32'h431b5986, 32'hc21784ba} /* (17, 10, 24) {real, imag} */,
  {32'hc22d593c, 32'hc132da34} /* (17, 10, 23) {real, imag} */,
  {32'hc1a043d6, 32'h414bed90} /* (17, 10, 22) {real, imag} */,
  {32'hc0c6cad0, 32'h4252033b} /* (17, 10, 21) {real, imag} */,
  {32'hc2b09d6e, 32'h422cc130} /* (17, 10, 20) {real, imag} */,
  {32'h42214e05, 32'h42d6a1b4} /* (17, 10, 19) {real, imag} */,
  {32'hc28a42d9, 32'h422897be} /* (17, 10, 18) {real, imag} */,
  {32'hc205b654, 32'h41fbaba2} /* (17, 10, 17) {real, imag} */,
  {32'hc1f125fa, 32'h00000000} /* (17, 10, 16) {real, imag} */,
  {32'hc205b654, 32'hc1fbaba2} /* (17, 10, 15) {real, imag} */,
  {32'hc28a42d9, 32'hc22897be} /* (17, 10, 14) {real, imag} */,
  {32'h42214e05, 32'hc2d6a1b4} /* (17, 10, 13) {real, imag} */,
  {32'hc2b09d6e, 32'hc22cc130} /* (17, 10, 12) {real, imag} */,
  {32'hc0c6cad0, 32'hc252033b} /* (17, 10, 11) {real, imag} */,
  {32'hc1a043d6, 32'hc14bed90} /* (17, 10, 10) {real, imag} */,
  {32'hc22d593c, 32'h4132da34} /* (17, 10, 9) {real, imag} */,
  {32'h431b5986, 32'h421784ba} /* (17, 10, 8) {real, imag} */,
  {32'h42097e23, 32'hc0925464} /* (17, 10, 7) {real, imag} */,
  {32'h42576b46, 32'h4095d880} /* (17, 10, 6) {real, imag} */,
  {32'h420b9c1c, 32'h408e2390} /* (17, 10, 5) {real, imag} */,
  {32'hc2c86064, 32'h42ac9e55} /* (17, 10, 4) {real, imag} */,
  {32'h42a5acdc, 32'hc2f3c40e} /* (17, 10, 3) {real, imag} */,
  {32'h42a17488, 32'h42281cdd} /* (17, 10, 2) {real, imag} */,
  {32'hc42abf33, 32'hc404f355} /* (17, 10, 1) {real, imag} */,
  {32'hc3876446, 32'h00000000} /* (17, 10, 0) {real, imag} */,
  {32'hc4c1ac54, 32'h44146a28} /* (17, 9, 31) {real, imag} */,
  {32'h4409e449, 32'hc31f7fa8} /* (17, 9, 30) {real, imag} */,
  {32'hc2e425ac, 32'h42ea709e} /* (17, 9, 29) {real, imag} */,
  {32'h4113f150, 32'h419fb9aa} /* (17, 9, 28) {real, imag} */,
  {32'h41ba7e68, 32'h41107768} /* (17, 9, 27) {real, imag} */,
  {32'hc2f58972, 32'hc1948a80} /* (17, 9, 26) {real, imag} */,
  {32'hc1c0cda2, 32'h42bb240c} /* (17, 9, 25) {real, imag} */,
  {32'h42798ac2, 32'hc2a1af17} /* (17, 9, 24) {real, imag} */,
  {32'hc0f8f8b0, 32'hc20eac36} /* (17, 9, 23) {real, imag} */,
  {32'h42573d8b, 32'h41aebb65} /* (17, 9, 22) {real, imag} */,
  {32'h42a1a650, 32'hc2cb45c0} /* (17, 9, 21) {real, imag} */,
  {32'hc27e28b9, 32'h4022a71c} /* (17, 9, 20) {real, imag} */,
  {32'hc12da776, 32'h424c529a} /* (17, 9, 19) {real, imag} */,
  {32'hbeac4540, 32'hc2997b07} /* (17, 9, 18) {real, imag} */,
  {32'h411d10d2, 32'hc2954d4c} /* (17, 9, 17) {real, imag} */,
  {32'h40f6110c, 32'h00000000} /* (17, 9, 16) {real, imag} */,
  {32'h411d10d2, 32'h42954d4c} /* (17, 9, 15) {real, imag} */,
  {32'hbeac4540, 32'h42997b07} /* (17, 9, 14) {real, imag} */,
  {32'hc12da776, 32'hc24c529a} /* (17, 9, 13) {real, imag} */,
  {32'hc27e28b9, 32'hc022a71c} /* (17, 9, 12) {real, imag} */,
  {32'h42a1a650, 32'h42cb45c0} /* (17, 9, 11) {real, imag} */,
  {32'h42573d8b, 32'hc1aebb65} /* (17, 9, 10) {real, imag} */,
  {32'hc0f8f8b0, 32'h420eac36} /* (17, 9, 9) {real, imag} */,
  {32'h42798ac2, 32'h42a1af17} /* (17, 9, 8) {real, imag} */,
  {32'hc1c0cda2, 32'hc2bb240c} /* (17, 9, 7) {real, imag} */,
  {32'hc2f58972, 32'h41948a80} /* (17, 9, 6) {real, imag} */,
  {32'h41ba7e68, 32'hc1107768} /* (17, 9, 5) {real, imag} */,
  {32'h4113f150, 32'hc19fb9aa} /* (17, 9, 4) {real, imag} */,
  {32'hc2e425ac, 32'hc2ea709e} /* (17, 9, 3) {real, imag} */,
  {32'h4409e449, 32'h431f7fa8} /* (17, 9, 2) {real, imag} */,
  {32'hc4c1ac54, 32'hc4146a28} /* (17, 9, 1) {real, imag} */,
  {32'hc4716984, 32'h00000000} /* (17, 9, 0) {real, imag} */,
  {32'hc501ec33, 32'h4439d1de} /* (17, 8, 31) {real, imag} */,
  {32'h442a9b16, 32'hc389b6ce} /* (17, 8, 30) {real, imag} */,
  {32'hc2dac762, 32'h42b32741} /* (17, 8, 29) {real, imag} */,
  {32'h421e9cf0, 32'hc2aa3fdd} /* (17, 8, 28) {real, imag} */,
  {32'h4255e068, 32'h4130e9b8} /* (17, 8, 27) {real, imag} */,
  {32'hc207fd9c, 32'h42e208fc} /* (17, 8, 26) {real, imag} */,
  {32'hc323766c, 32'h427d7860} /* (17, 8, 25) {real, imag} */,
  {32'h429d3498, 32'hc2466197} /* (17, 8, 24) {real, imag} */,
  {32'hc1ace50d, 32'hc20887bc} /* (17, 8, 23) {real, imag} */,
  {32'h43220ca4, 32'hc29c2a35} /* (17, 8, 22) {real, imag} */,
  {32'h42034afa, 32'h42b1bf94} /* (17, 8, 21) {real, imag} */,
  {32'h428fb01b, 32'h4115e1c8} /* (17, 8, 20) {real, imag} */,
  {32'hc1e4111c, 32'hc2194b44} /* (17, 8, 19) {real, imag} */,
  {32'h4187a5f4, 32'h417d0070} /* (17, 8, 18) {real, imag} */,
  {32'hc2ba7651, 32'hc1aff336} /* (17, 8, 17) {real, imag} */,
  {32'h425d4780, 32'h00000000} /* (17, 8, 16) {real, imag} */,
  {32'hc2ba7651, 32'h41aff336} /* (17, 8, 15) {real, imag} */,
  {32'h4187a5f4, 32'hc17d0070} /* (17, 8, 14) {real, imag} */,
  {32'hc1e4111c, 32'h42194b44} /* (17, 8, 13) {real, imag} */,
  {32'h428fb01b, 32'hc115e1c8} /* (17, 8, 12) {real, imag} */,
  {32'h42034afa, 32'hc2b1bf94} /* (17, 8, 11) {real, imag} */,
  {32'h43220ca4, 32'h429c2a35} /* (17, 8, 10) {real, imag} */,
  {32'hc1ace50d, 32'h420887bc} /* (17, 8, 9) {real, imag} */,
  {32'h429d3498, 32'h42466197} /* (17, 8, 8) {real, imag} */,
  {32'hc323766c, 32'hc27d7860} /* (17, 8, 7) {real, imag} */,
  {32'hc207fd9c, 32'hc2e208fc} /* (17, 8, 6) {real, imag} */,
  {32'h4255e068, 32'hc130e9b8} /* (17, 8, 5) {real, imag} */,
  {32'h421e9cf0, 32'h42aa3fdd} /* (17, 8, 4) {real, imag} */,
  {32'hc2dac762, 32'hc2b32741} /* (17, 8, 3) {real, imag} */,
  {32'h442a9b16, 32'h4389b6ce} /* (17, 8, 2) {real, imag} */,
  {32'hc501ec33, 32'hc439d1de} /* (17, 8, 1) {real, imag} */,
  {32'hc4c992a0, 32'h00000000} /* (17, 8, 0) {real, imag} */,
  {32'hc511af73, 32'h447b6594} /* (17, 7, 31) {real, imag} */,
  {32'h44265415, 32'hc3c11770} /* (17, 7, 30) {real, imag} */,
  {32'hc275c959, 32'h426fe26a} /* (17, 7, 29) {real, imag} */,
  {32'hc2d68f79, 32'h42fcdeb2} /* (17, 7, 28) {real, imag} */,
  {32'h43624e79, 32'hc2bf5c15} /* (17, 7, 27) {real, imag} */,
  {32'h41aa2fea, 32'h43332cde} /* (17, 7, 26) {real, imag} */,
  {32'hc237d7bc, 32'hc0327200} /* (17, 7, 25) {real, imag} */,
  {32'h42e30000, 32'hc19faf70} /* (17, 7, 24) {real, imag} */,
  {32'h431cf546, 32'h41cacbda} /* (17, 7, 23) {real, imag} */,
  {32'hc23ec6d5, 32'hc287f47a} /* (17, 7, 22) {real, imag} */,
  {32'hc1aa9380, 32'h422f33a2} /* (17, 7, 21) {real, imag} */,
  {32'h41b7fb5a, 32'h41d39ca2} /* (17, 7, 20) {real, imag} */,
  {32'h4205a654, 32'hc2877c39} /* (17, 7, 19) {real, imag} */,
  {32'h42478d77, 32'hc0903d30} /* (17, 7, 18) {real, imag} */,
  {32'hc0ed25e9, 32'h42a575e5} /* (17, 7, 17) {real, imag} */,
  {32'h42c1c11c, 32'h00000000} /* (17, 7, 16) {real, imag} */,
  {32'hc0ed25e9, 32'hc2a575e5} /* (17, 7, 15) {real, imag} */,
  {32'h42478d77, 32'h40903d30} /* (17, 7, 14) {real, imag} */,
  {32'h4205a654, 32'h42877c39} /* (17, 7, 13) {real, imag} */,
  {32'h41b7fb5a, 32'hc1d39ca2} /* (17, 7, 12) {real, imag} */,
  {32'hc1aa9380, 32'hc22f33a2} /* (17, 7, 11) {real, imag} */,
  {32'hc23ec6d5, 32'h4287f47a} /* (17, 7, 10) {real, imag} */,
  {32'h431cf546, 32'hc1cacbda} /* (17, 7, 9) {real, imag} */,
  {32'h42e30000, 32'h419faf70} /* (17, 7, 8) {real, imag} */,
  {32'hc237d7bc, 32'h40327200} /* (17, 7, 7) {real, imag} */,
  {32'h41aa2fea, 32'hc3332cde} /* (17, 7, 6) {real, imag} */,
  {32'h43624e79, 32'h42bf5c15} /* (17, 7, 5) {real, imag} */,
  {32'hc2d68f79, 32'hc2fcdeb2} /* (17, 7, 4) {real, imag} */,
  {32'hc275c959, 32'hc26fe26a} /* (17, 7, 3) {real, imag} */,
  {32'h44265415, 32'h43c11770} /* (17, 7, 2) {real, imag} */,
  {32'hc511af73, 32'hc47b6594} /* (17, 7, 1) {real, imag} */,
  {32'hc50588ca, 32'h00000000} /* (17, 7, 0) {real, imag} */,
  {32'hc51250b1, 32'h449bcfa8} /* (17, 6, 31) {real, imag} */,
  {32'h441716c9, 32'hc3d22a1e} /* (17, 6, 30) {real, imag} */,
  {32'hc2c2013a, 32'h419308cb} /* (17, 6, 29) {real, imag} */,
  {32'hc2b0bf4a, 32'h42405354} /* (17, 6, 28) {real, imag} */,
  {32'h437bbe72, 32'h410f35c2} /* (17, 6, 27) {real, imag} */,
  {32'h4307894c, 32'h42cf6074} /* (17, 6, 26) {real, imag} */,
  {32'h40513f98, 32'h418668f3} /* (17, 6, 25) {real, imag} */,
  {32'h42397fde, 32'hc32ccfe1} /* (17, 6, 24) {real, imag} */,
  {32'hc1af5e02, 32'h42227b78} /* (17, 6, 23) {real, imag} */,
  {32'h40d9e1e2, 32'h4265288e} /* (17, 6, 22) {real, imag} */,
  {32'hc1a05fda, 32'hc31d1f4d} /* (17, 6, 21) {real, imag} */,
  {32'hc0e0d79c, 32'hc266b78a} /* (17, 6, 20) {real, imag} */,
  {32'h42cea7da, 32'h424c9b5c} /* (17, 6, 19) {real, imag} */,
  {32'hbecdd580, 32'h40bd7b3c} /* (17, 6, 18) {real, imag} */,
  {32'hc22d5138, 32'h3e30eb80} /* (17, 6, 17) {real, imag} */,
  {32'h4165e090, 32'h00000000} /* (17, 6, 16) {real, imag} */,
  {32'hc22d5138, 32'hbe30eb80} /* (17, 6, 15) {real, imag} */,
  {32'hbecdd580, 32'hc0bd7b3c} /* (17, 6, 14) {real, imag} */,
  {32'h42cea7da, 32'hc24c9b5c} /* (17, 6, 13) {real, imag} */,
  {32'hc0e0d79c, 32'h4266b78a} /* (17, 6, 12) {real, imag} */,
  {32'hc1a05fda, 32'h431d1f4d} /* (17, 6, 11) {real, imag} */,
  {32'h40d9e1e2, 32'hc265288e} /* (17, 6, 10) {real, imag} */,
  {32'hc1af5e02, 32'hc2227b78} /* (17, 6, 9) {real, imag} */,
  {32'h42397fde, 32'h432ccfe1} /* (17, 6, 8) {real, imag} */,
  {32'h40513f98, 32'hc18668f3} /* (17, 6, 7) {real, imag} */,
  {32'h4307894c, 32'hc2cf6074} /* (17, 6, 6) {real, imag} */,
  {32'h437bbe72, 32'hc10f35c2} /* (17, 6, 5) {real, imag} */,
  {32'hc2b0bf4a, 32'hc2405354} /* (17, 6, 4) {real, imag} */,
  {32'hc2c2013a, 32'hc19308cb} /* (17, 6, 3) {real, imag} */,
  {32'h441716c9, 32'h43d22a1e} /* (17, 6, 2) {real, imag} */,
  {32'hc51250b1, 32'hc49bcfa8} /* (17, 6, 1) {real, imag} */,
  {32'hc5139320, 32'h00000000} /* (17, 6, 0) {real, imag} */,
  {32'hc4fb552a, 32'h44d553d6} /* (17, 5, 31) {real, imag} */,
  {32'h42e1bf04, 32'hc4201d84} /* (17, 5, 30) {real, imag} */,
  {32'hc22352c8, 32'h422e8af0} /* (17, 5, 29) {real, imag} */,
  {32'h4328a59d, 32'hc13b53b0} /* (17, 5, 28) {real, imag} */,
  {32'h42e9cc16, 32'h422b1b84} /* (17, 5, 27) {real, imag} */,
  {32'h429d635b, 32'h42ce357b} /* (17, 5, 26) {real, imag} */,
  {32'h423b2a19, 32'hc24703ea} /* (17, 5, 25) {real, imag} */,
  {32'hc2a65265, 32'hc2ed30c9} /* (17, 5, 24) {real, imag} */,
  {32'hc11d1530, 32'hc136c06c} /* (17, 5, 23) {real, imag} */,
  {32'hc0f35020, 32'h42b72697} /* (17, 5, 22) {real, imag} */,
  {32'h42881374, 32'hc25b4cfa} /* (17, 5, 21) {real, imag} */,
  {32'h40822628, 32'h411f79ea} /* (17, 5, 20) {real, imag} */,
  {32'hc225c5e9, 32'h428ae2d6} /* (17, 5, 19) {real, imag} */,
  {32'hc2152024, 32'h4220ec48} /* (17, 5, 18) {real, imag} */,
  {32'h4156a7dd, 32'h424a653a} /* (17, 5, 17) {real, imag} */,
  {32'hc212c157, 32'h00000000} /* (17, 5, 16) {real, imag} */,
  {32'h4156a7dd, 32'hc24a653a} /* (17, 5, 15) {real, imag} */,
  {32'hc2152024, 32'hc220ec48} /* (17, 5, 14) {real, imag} */,
  {32'hc225c5e9, 32'hc28ae2d6} /* (17, 5, 13) {real, imag} */,
  {32'h40822628, 32'hc11f79ea} /* (17, 5, 12) {real, imag} */,
  {32'h42881374, 32'h425b4cfa} /* (17, 5, 11) {real, imag} */,
  {32'hc0f35020, 32'hc2b72697} /* (17, 5, 10) {real, imag} */,
  {32'hc11d1530, 32'h4136c06c} /* (17, 5, 9) {real, imag} */,
  {32'hc2a65265, 32'h42ed30c9} /* (17, 5, 8) {real, imag} */,
  {32'h423b2a19, 32'h424703ea} /* (17, 5, 7) {real, imag} */,
  {32'h429d635b, 32'hc2ce357b} /* (17, 5, 6) {real, imag} */,
  {32'h42e9cc16, 32'hc22b1b84} /* (17, 5, 5) {real, imag} */,
  {32'h4328a59d, 32'h413b53b0} /* (17, 5, 4) {real, imag} */,
  {32'hc22352c8, 32'hc22e8af0} /* (17, 5, 3) {real, imag} */,
  {32'h42e1bf04, 32'h44201d84} /* (17, 5, 2) {real, imag} */,
  {32'hc4fb552a, 32'hc4d553d6} /* (17, 5, 1) {real, imag} */,
  {32'hc51cb4bc, 32'h00000000} /* (17, 5, 0) {real, imag} */,
  {32'hc4dab882, 32'h44fff7d5} /* (17, 4, 31) {real, imag} */,
  {32'hc3936a08, 32'hc43dcaf5} /* (17, 4, 30) {real, imag} */,
  {32'h421f6f0e, 32'h413f044a} /* (17, 4, 29) {real, imag} */,
  {32'h438675be, 32'hc27659f0} /* (17, 4, 28) {real, imag} */,
  {32'h4357a466, 32'h4350191b} /* (17, 4, 27) {real, imag} */,
  {32'hc2c347c8, 32'h417b7e1a} /* (17, 4, 26) {real, imag} */,
  {32'h4217e6b3, 32'h42064b8b} /* (17, 4, 25) {real, imag} */,
  {32'hc2a9fc7e, 32'hc2bf31ef} /* (17, 4, 24) {real, imag} */,
  {32'h424b83fb, 32'h3fe2fbb0} /* (17, 4, 23) {real, imag} */,
  {32'hc24a0ff2, 32'hc2a953e1} /* (17, 4, 22) {real, imag} */,
  {32'hbffaabf0, 32'hc2380f8f} /* (17, 4, 21) {real, imag} */,
  {32'h42e8a025, 32'hc1a96e1a} /* (17, 4, 20) {real, imag} */,
  {32'hc1e62fe8, 32'h420fac7a} /* (17, 4, 19) {real, imag} */,
  {32'h414df0e0, 32'hc08681f0} /* (17, 4, 18) {real, imag} */,
  {32'hc2886e92, 32'h427a7ad2} /* (17, 4, 17) {real, imag} */,
  {32'h4249ba34, 32'h00000000} /* (17, 4, 16) {real, imag} */,
  {32'hc2886e92, 32'hc27a7ad2} /* (17, 4, 15) {real, imag} */,
  {32'h414df0e0, 32'h408681f0} /* (17, 4, 14) {real, imag} */,
  {32'hc1e62fe8, 32'hc20fac7a} /* (17, 4, 13) {real, imag} */,
  {32'h42e8a025, 32'h41a96e1a} /* (17, 4, 12) {real, imag} */,
  {32'hbffaabf0, 32'h42380f8f} /* (17, 4, 11) {real, imag} */,
  {32'hc24a0ff2, 32'h42a953e1} /* (17, 4, 10) {real, imag} */,
  {32'h424b83fb, 32'hbfe2fbb0} /* (17, 4, 9) {real, imag} */,
  {32'hc2a9fc7e, 32'h42bf31ef} /* (17, 4, 8) {real, imag} */,
  {32'h4217e6b3, 32'hc2064b8b} /* (17, 4, 7) {real, imag} */,
  {32'hc2c347c8, 32'hc17b7e1a} /* (17, 4, 6) {real, imag} */,
  {32'h4357a466, 32'hc350191b} /* (17, 4, 5) {real, imag} */,
  {32'h438675be, 32'h427659f0} /* (17, 4, 4) {real, imag} */,
  {32'h421f6f0e, 32'hc13f044a} /* (17, 4, 3) {real, imag} */,
  {32'hc3936a08, 32'h443dcaf5} /* (17, 4, 2) {real, imag} */,
  {32'hc4dab882, 32'hc4fff7d5} /* (17, 4, 1) {real, imag} */,
  {32'hc5158ece, 32'h00000000} /* (17, 4, 0) {real, imag} */,
  {32'hc4e0f38d, 32'h4511965f} /* (17, 3, 31) {real, imag} */,
  {32'hc3ad3484, 32'hc4718cae} /* (17, 3, 30) {real, imag} */,
  {32'h43512bb7, 32'h433a35be} /* (17, 3, 29) {real, imag} */,
  {32'h434ce992, 32'hc31374fc} /* (17, 3, 28) {real, imag} */,
  {32'h43187c8c, 32'h43988bda} /* (17, 3, 27) {real, imag} */,
  {32'h4223331c, 32'hc297d7cc} /* (17, 3, 26) {real, imag} */,
  {32'hc0c77178, 32'h428bdf7c} /* (17, 3, 25) {real, imag} */,
  {32'h4290761d, 32'hc2fff03a} /* (17, 3, 24) {real, imag} */,
  {32'hbf53b6c0, 32'hc22bc019} /* (17, 3, 23) {real, imag} */,
  {32'h4012bb30, 32'hc297c268} /* (17, 3, 22) {real, imag} */,
  {32'h418fac80, 32'hc3237b58} /* (17, 3, 21) {real, imag} */,
  {32'hc1aa46b8, 32'h4140cacf} /* (17, 3, 20) {real, imag} */,
  {32'hc1cdf184, 32'h416c31aa} /* (17, 3, 19) {real, imag} */,
  {32'hc2f5c0ca, 32'h413e3965} /* (17, 3, 18) {real, imag} */,
  {32'h4282d3e1, 32'hc1c47176} /* (17, 3, 17) {real, imag} */,
  {32'hc297cee8, 32'h00000000} /* (17, 3, 16) {real, imag} */,
  {32'h4282d3e1, 32'h41c47176} /* (17, 3, 15) {real, imag} */,
  {32'hc2f5c0ca, 32'hc13e3965} /* (17, 3, 14) {real, imag} */,
  {32'hc1cdf184, 32'hc16c31aa} /* (17, 3, 13) {real, imag} */,
  {32'hc1aa46b8, 32'hc140cacf} /* (17, 3, 12) {real, imag} */,
  {32'h418fac80, 32'h43237b58} /* (17, 3, 11) {real, imag} */,
  {32'h4012bb30, 32'h4297c268} /* (17, 3, 10) {real, imag} */,
  {32'hbf53b6c0, 32'h422bc019} /* (17, 3, 9) {real, imag} */,
  {32'h4290761d, 32'h42fff03a} /* (17, 3, 8) {real, imag} */,
  {32'hc0c77178, 32'hc28bdf7c} /* (17, 3, 7) {real, imag} */,
  {32'h4223331c, 32'h4297d7cc} /* (17, 3, 6) {real, imag} */,
  {32'h43187c8c, 32'hc3988bda} /* (17, 3, 5) {real, imag} */,
  {32'h434ce992, 32'h431374fc} /* (17, 3, 4) {real, imag} */,
  {32'h43512bb7, 32'hc33a35be} /* (17, 3, 3) {real, imag} */,
  {32'hc3ad3484, 32'h44718cae} /* (17, 3, 2) {real, imag} */,
  {32'hc4e0f38d, 32'hc511965f} /* (17, 3, 1) {real, imag} */,
  {32'hc513893a, 32'h00000000} /* (17, 3, 0) {real, imag} */,
  {32'hc4d14def, 32'h45071064} /* (17, 2, 31) {real, imag} */,
  {32'hc3b35f0e, 32'hc471e9ba} /* (17, 2, 30) {real, imag} */,
  {32'h43937a69, 32'h43748ee4} /* (17, 2, 29) {real, imag} */,
  {32'h417a4100, 32'hc3b8ec6c} /* (17, 2, 28) {real, imag} */,
  {32'h429ecc7e, 32'h43791de1} /* (17, 2, 27) {real, imag} */,
  {32'h427cbdb9, 32'hc2c81c10} /* (17, 2, 26) {real, imag} */,
  {32'hc28607b5, 32'h430f4e9f} /* (17, 2, 25) {real, imag} */,
  {32'h42f93f04, 32'hc3199ea5} /* (17, 2, 24) {real, imag} */,
  {32'hc264bb9c, 32'hc2945600} /* (17, 2, 23) {real, imag} */,
  {32'h4217098d, 32'hc1b03a46} /* (17, 2, 22) {real, imag} */,
  {32'hc2bc9ef6, 32'hc2bbe582} /* (17, 2, 21) {real, imag} */,
  {32'h429f080e, 32'h42aca09e} /* (17, 2, 20) {real, imag} */,
  {32'hc1c9237e, 32'h4239a0ec} /* (17, 2, 19) {real, imag} */,
  {32'hc1e6254e, 32'hc2113a52} /* (17, 2, 18) {real, imag} */,
  {32'h42a8071e, 32'h415efe90} /* (17, 2, 17) {real, imag} */,
  {32'hc2faf381, 32'h00000000} /* (17, 2, 16) {real, imag} */,
  {32'h42a8071e, 32'hc15efe90} /* (17, 2, 15) {real, imag} */,
  {32'hc1e6254e, 32'h42113a52} /* (17, 2, 14) {real, imag} */,
  {32'hc1c9237e, 32'hc239a0ec} /* (17, 2, 13) {real, imag} */,
  {32'h429f080e, 32'hc2aca09e} /* (17, 2, 12) {real, imag} */,
  {32'hc2bc9ef6, 32'h42bbe582} /* (17, 2, 11) {real, imag} */,
  {32'h4217098d, 32'h41b03a46} /* (17, 2, 10) {real, imag} */,
  {32'hc264bb9c, 32'h42945600} /* (17, 2, 9) {real, imag} */,
  {32'h42f93f04, 32'h43199ea5} /* (17, 2, 8) {real, imag} */,
  {32'hc28607b5, 32'hc30f4e9f} /* (17, 2, 7) {real, imag} */,
  {32'h427cbdb9, 32'h42c81c10} /* (17, 2, 6) {real, imag} */,
  {32'h429ecc7e, 32'hc3791de1} /* (17, 2, 5) {real, imag} */,
  {32'h417a4100, 32'h43b8ec6c} /* (17, 2, 4) {real, imag} */,
  {32'h43937a69, 32'hc3748ee4} /* (17, 2, 3) {real, imag} */,
  {32'hc3b35f0e, 32'h4471e9ba} /* (17, 2, 2) {real, imag} */,
  {32'hc4d14def, 32'hc5071064} /* (17, 2, 1) {real, imag} */,
  {32'hc51b9977, 32'h00000000} /* (17, 2, 0) {real, imag} */,
  {32'hc4d0e884, 32'h44f913cb} /* (17, 1, 31) {real, imag} */,
  {32'hc341b94a, 32'hc461c57b} /* (17, 1, 30) {real, imag} */,
  {32'h4360b47e, 32'h4361d376} /* (17, 1, 29) {real, imag} */,
  {32'h41eafe4c, 32'hc3be165d} /* (17, 1, 28) {real, imag} */,
  {32'h42fb813f, 32'h4378ffef} /* (17, 1, 27) {real, imag} */,
  {32'hc224a1f1, 32'hc29e9be4} /* (17, 1, 26) {real, imag} */,
  {32'hc2369183, 32'h429eda2a} /* (17, 1, 25) {real, imag} */,
  {32'h419a73ad, 32'hc2f4b0d2} /* (17, 1, 24) {real, imag} */,
  {32'h4160e0d2, 32'hc2d4fb20} /* (17, 1, 23) {real, imag} */,
  {32'hc0aebf30, 32'hc20113c5} /* (17, 1, 22) {real, imag} */,
  {32'h419bec44, 32'hc1c197b6} /* (17, 1, 21) {real, imag} */,
  {32'h42ab70e6, 32'h4231136e} /* (17, 1, 20) {real, imag} */,
  {32'hc1131816, 32'hc1aabd5c} /* (17, 1, 19) {real, imag} */,
  {32'hc1ca334b, 32'h42c5c9fe} /* (17, 1, 18) {real, imag} */,
  {32'h41efdf1f, 32'hc1a4dca3} /* (17, 1, 17) {real, imag} */,
  {32'h41d73a1d, 32'h00000000} /* (17, 1, 16) {real, imag} */,
  {32'h41efdf1f, 32'h41a4dca3} /* (17, 1, 15) {real, imag} */,
  {32'hc1ca334b, 32'hc2c5c9fe} /* (17, 1, 14) {real, imag} */,
  {32'hc1131816, 32'h41aabd5c} /* (17, 1, 13) {real, imag} */,
  {32'h42ab70e6, 32'hc231136e} /* (17, 1, 12) {real, imag} */,
  {32'h419bec44, 32'h41c197b6} /* (17, 1, 11) {real, imag} */,
  {32'hc0aebf30, 32'h420113c5} /* (17, 1, 10) {real, imag} */,
  {32'h4160e0d2, 32'h42d4fb20} /* (17, 1, 9) {real, imag} */,
  {32'h419a73ad, 32'h42f4b0d2} /* (17, 1, 8) {real, imag} */,
  {32'hc2369183, 32'hc29eda2a} /* (17, 1, 7) {real, imag} */,
  {32'hc224a1f1, 32'h429e9be4} /* (17, 1, 6) {real, imag} */,
  {32'h42fb813f, 32'hc378ffef} /* (17, 1, 5) {real, imag} */,
  {32'h41eafe4c, 32'h43be165d} /* (17, 1, 4) {real, imag} */,
  {32'h4360b47e, 32'hc361d376} /* (17, 1, 3) {real, imag} */,
  {32'hc341b94a, 32'h4461c57b} /* (17, 1, 2) {real, imag} */,
  {32'hc4d0e884, 32'hc4f913cb} /* (17, 1, 1) {real, imag} */,
  {32'hc528b830, 32'h00000000} /* (17, 1, 0) {real, imag} */,
  {32'hc4dfa87c, 32'h44c76120} /* (17, 0, 31) {real, imag} */,
  {32'h42625df0, 32'hc41ba575} /* (17, 0, 30) {real, imag} */,
  {32'h42baf1f5, 32'h430110fc} /* (17, 0, 29) {real, imag} */,
  {32'h4142cf00, 32'hc2d01c08} /* (17, 0, 28) {real, imag} */,
  {32'h4294237f, 32'hc126b8a8} /* (17, 0, 27) {real, imag} */,
  {32'h41e6fb1b, 32'h3e85f680} /* (17, 0, 26) {real, imag} */,
  {32'hc19e17c8, 32'h428427ae} /* (17, 0, 25) {real, imag} */,
  {32'h42096f4e, 32'hc1036f94} /* (17, 0, 24) {real, imag} */,
  {32'h41c69ab2, 32'h413fe33c} /* (17, 0, 23) {real, imag} */,
  {32'hc208d186, 32'h4188848d} /* (17, 0, 22) {real, imag} */,
  {32'hc18f24c2, 32'h41c571a4} /* (17, 0, 21) {real, imag} */,
  {32'h42283c5c, 32'h423c3370} /* (17, 0, 20) {real, imag} */,
  {32'hc16396c1, 32'h41f4d766} /* (17, 0, 19) {real, imag} */,
  {32'h415158d8, 32'h42071ebe} /* (17, 0, 18) {real, imag} */,
  {32'hc159425c, 32'h3fa80050} /* (17, 0, 17) {real, imag} */,
  {32'h41627f9c, 32'h00000000} /* (17, 0, 16) {real, imag} */,
  {32'hc159425c, 32'hbfa80050} /* (17, 0, 15) {real, imag} */,
  {32'h415158d8, 32'hc2071ebe} /* (17, 0, 14) {real, imag} */,
  {32'hc16396c1, 32'hc1f4d766} /* (17, 0, 13) {real, imag} */,
  {32'h42283c5c, 32'hc23c3370} /* (17, 0, 12) {real, imag} */,
  {32'hc18f24c2, 32'hc1c571a4} /* (17, 0, 11) {real, imag} */,
  {32'hc208d186, 32'hc188848d} /* (17, 0, 10) {real, imag} */,
  {32'h41c69ab2, 32'hc13fe33c} /* (17, 0, 9) {real, imag} */,
  {32'h42096f4e, 32'h41036f94} /* (17, 0, 8) {real, imag} */,
  {32'hc19e17c8, 32'hc28427ae} /* (17, 0, 7) {real, imag} */,
  {32'h41e6fb1b, 32'hbe85f680} /* (17, 0, 6) {real, imag} */,
  {32'h4294237f, 32'h4126b8a8} /* (17, 0, 5) {real, imag} */,
  {32'h4142cf00, 32'h42d01c08} /* (17, 0, 4) {real, imag} */,
  {32'h42baf1f5, 32'hc30110fc} /* (17, 0, 3) {real, imag} */,
  {32'h42625df0, 32'h441ba575} /* (17, 0, 2) {real, imag} */,
  {32'hc4dfa87c, 32'hc4c76120} /* (17, 0, 1) {real, imag} */,
  {32'hc51fc958, 32'h00000000} /* (17, 0, 0) {real, imag} */,
  {32'hc44cda95, 32'h439cadae} /* (16, 31, 31) {real, imag} */,
  {32'h432d539a, 32'hc37c54be} /* (16, 31, 30) {real, imag} */,
  {32'h424da90e, 32'h42a4fe42} /* (16, 31, 29) {real, imag} */,
  {32'hc29b9a69, 32'h42795a4e} /* (16, 31, 28) {real, imag} */,
  {32'h42d4e3ad, 32'hc1c4dff0} /* (16, 31, 27) {real, imag} */,
  {32'h4221b926, 32'hc1544bd4} /* (16, 31, 26) {real, imag} */,
  {32'hc1aed732, 32'h40589470} /* (16, 31, 25) {real, imag} */,
  {32'h40129328, 32'h4289d4c5} /* (16, 31, 24) {real, imag} */,
  {32'hc1488120, 32'hc14e57c5} /* (16, 31, 23) {real, imag} */,
  {32'h40523fdc, 32'hc0188e58} /* (16, 31, 22) {real, imag} */,
  {32'h41554c0a, 32'h41fcd610} /* (16, 31, 21) {real, imag} */,
  {32'hc086c5fe, 32'h40a12d20} /* (16, 31, 20) {real, imag} */,
  {32'hc2c628ac, 32'hc2b52652} /* (16, 31, 19) {real, imag} */,
  {32'h422d493a, 32'hc2211fe3} /* (16, 31, 18) {real, imag} */,
  {32'h416efa24, 32'hc1abedb0} /* (16, 31, 17) {real, imag} */,
  {32'h42ab895e, 32'h00000000} /* (16, 31, 16) {real, imag} */,
  {32'h416efa24, 32'h41abedb0} /* (16, 31, 15) {real, imag} */,
  {32'h422d493a, 32'h42211fe3} /* (16, 31, 14) {real, imag} */,
  {32'hc2c628ac, 32'h42b52652} /* (16, 31, 13) {real, imag} */,
  {32'hc086c5fe, 32'hc0a12d20} /* (16, 31, 12) {real, imag} */,
  {32'h41554c0a, 32'hc1fcd610} /* (16, 31, 11) {real, imag} */,
  {32'h40523fdc, 32'h40188e58} /* (16, 31, 10) {real, imag} */,
  {32'hc1488120, 32'h414e57c5} /* (16, 31, 9) {real, imag} */,
  {32'h40129328, 32'hc289d4c5} /* (16, 31, 8) {real, imag} */,
  {32'hc1aed732, 32'hc0589470} /* (16, 31, 7) {real, imag} */,
  {32'h4221b926, 32'h41544bd4} /* (16, 31, 6) {real, imag} */,
  {32'h42d4e3ad, 32'h41c4dff0} /* (16, 31, 5) {real, imag} */,
  {32'hc29b9a69, 32'hc2795a4e} /* (16, 31, 4) {real, imag} */,
  {32'h424da90e, 32'hc2a4fe42} /* (16, 31, 3) {real, imag} */,
  {32'h432d539a, 32'h437c54be} /* (16, 31, 2) {real, imag} */,
  {32'hc44cda95, 32'hc39cadae} /* (16, 31, 1) {real, imag} */,
  {32'hc48fd602, 32'h00000000} /* (16, 31, 0) {real, imag} */,
  {32'hc495eedc, 32'h43168e68} /* (16, 30, 31) {real, imag} */,
  {32'h43a675da, 32'hc327c75e} /* (16, 30, 30) {real, imag} */,
  {32'h42d17991, 32'h42edc80e} /* (16, 30, 29) {real, imag} */,
  {32'hc1d8ec1d, 32'h41c33e10} /* (16, 30, 28) {real, imag} */,
  {32'h4347428f, 32'hc2ef2d26} /* (16, 30, 27) {real, imag} */,
  {32'h42b82066, 32'hc2cdd6b0} /* (16, 30, 26) {real, imag} */,
  {32'hbfa6ff00, 32'h42fce8ee} /* (16, 30, 25) {real, imag} */,
  {32'hc1dd4c6e, 32'hbfa8e890} /* (16, 30, 24) {real, imag} */,
  {32'hbfc76180, 32'hc188bf60} /* (16, 30, 23) {real, imag} */,
  {32'hc182faa4, 32'hc222bac2} /* (16, 30, 22) {real, imag} */,
  {32'h4239959a, 32'hc1467b70} /* (16, 30, 21) {real, imag} */,
  {32'hc11b6472, 32'h41c3532d} /* (16, 30, 20) {real, imag} */,
  {32'hc21a6ca6, 32'h427d0f74} /* (16, 30, 19) {real, imag} */,
  {32'hc2a291f3, 32'h42a49903} /* (16, 30, 18) {real, imag} */,
  {32'hc1b2708a, 32'hc138b857} /* (16, 30, 17) {real, imag} */,
  {32'hc1879631, 32'h00000000} /* (16, 30, 16) {real, imag} */,
  {32'hc1b2708a, 32'h4138b857} /* (16, 30, 15) {real, imag} */,
  {32'hc2a291f3, 32'hc2a49903} /* (16, 30, 14) {real, imag} */,
  {32'hc21a6ca6, 32'hc27d0f74} /* (16, 30, 13) {real, imag} */,
  {32'hc11b6472, 32'hc1c3532d} /* (16, 30, 12) {real, imag} */,
  {32'h4239959a, 32'h41467b70} /* (16, 30, 11) {real, imag} */,
  {32'hc182faa4, 32'h4222bac2} /* (16, 30, 10) {real, imag} */,
  {32'hbfc76180, 32'h4188bf60} /* (16, 30, 9) {real, imag} */,
  {32'hc1dd4c6e, 32'h3fa8e890} /* (16, 30, 8) {real, imag} */,
  {32'hbfa6ff00, 32'hc2fce8ee} /* (16, 30, 7) {real, imag} */,
  {32'h42b82066, 32'h42cdd6b0} /* (16, 30, 6) {real, imag} */,
  {32'h4347428f, 32'h42ef2d26} /* (16, 30, 5) {real, imag} */,
  {32'hc1d8ec1d, 32'hc1c33e10} /* (16, 30, 4) {real, imag} */,
  {32'h42d17991, 32'hc2edc80e} /* (16, 30, 3) {real, imag} */,
  {32'h43a675da, 32'h4327c75e} /* (16, 30, 2) {real, imag} */,
  {32'hc495eedc, 32'hc3168e68} /* (16, 30, 1) {real, imag} */,
  {32'hc4908a20, 32'h00000000} /* (16, 30, 0) {real, imag} */,
  {32'hc4c948c1, 32'h42e088a4} /* (16, 29, 31) {real, imag} */,
  {32'h43d72d76, 32'hc3731e8a} /* (16, 29, 30) {real, imag} */,
  {32'h42a2dbdc, 32'h41939cdc} /* (16, 29, 29) {real, imag} */,
  {32'hc32578c0, 32'h40b4e0e0} /* (16, 29, 28) {real, imag} */,
  {32'h431b16f4, 32'hc3012303} /* (16, 29, 27) {real, imag} */,
  {32'h433a0d2e, 32'hc32f76af} /* (16, 29, 26) {real, imag} */,
  {32'hc27bd6f8, 32'hc21874b7} /* (16, 29, 25) {real, imag} */,
  {32'hc134f682, 32'h3f809300} /* (16, 29, 24) {real, imag} */,
  {32'h42c29442, 32'hc1326142} /* (16, 29, 23) {real, imag} */,
  {32'hc0948e22, 32'h4233c56a} /* (16, 29, 22) {real, imag} */,
  {32'hc1cd283c, 32'hc2856e87} /* (16, 29, 21) {real, imag} */,
  {32'hc24d840a, 32'h4122c8cc} /* (16, 29, 20) {real, imag} */,
  {32'h42913f64, 32'hc1b0156b} /* (16, 29, 19) {real, imag} */,
  {32'hc28e3966, 32'h422d200a} /* (16, 29, 18) {real, imag} */,
  {32'hc1589e56, 32'h42436710} /* (16, 29, 17) {real, imag} */,
  {32'hc1a61850, 32'h00000000} /* (16, 29, 16) {real, imag} */,
  {32'hc1589e56, 32'hc2436710} /* (16, 29, 15) {real, imag} */,
  {32'hc28e3966, 32'hc22d200a} /* (16, 29, 14) {real, imag} */,
  {32'h42913f64, 32'h41b0156b} /* (16, 29, 13) {real, imag} */,
  {32'hc24d840a, 32'hc122c8cc} /* (16, 29, 12) {real, imag} */,
  {32'hc1cd283c, 32'h42856e87} /* (16, 29, 11) {real, imag} */,
  {32'hc0948e22, 32'hc233c56a} /* (16, 29, 10) {real, imag} */,
  {32'h42c29442, 32'h41326142} /* (16, 29, 9) {real, imag} */,
  {32'hc134f682, 32'hbf809300} /* (16, 29, 8) {real, imag} */,
  {32'hc27bd6f8, 32'h421874b7} /* (16, 29, 7) {real, imag} */,
  {32'h433a0d2e, 32'h432f76af} /* (16, 29, 6) {real, imag} */,
  {32'h431b16f4, 32'h43012303} /* (16, 29, 5) {real, imag} */,
  {32'hc32578c0, 32'hc0b4e0e0} /* (16, 29, 4) {real, imag} */,
  {32'h42a2dbdc, 32'hc1939cdc} /* (16, 29, 3) {real, imag} */,
  {32'h43d72d76, 32'h43731e8a} /* (16, 29, 2) {real, imag} */,
  {32'hc4c948c1, 32'hc2e088a4} /* (16, 29, 1) {real, imag} */,
  {32'hc46a51fc, 32'h00000000} /* (16, 29, 0) {real, imag} */,
  {32'hc4ca6a6d, 32'h4335b078} /* (16, 28, 31) {real, imag} */,
  {32'h43dc085d, 32'hc39cced3} /* (16, 28, 30) {real, imag} */,
  {32'hc00235c8, 32'hc195f5be} /* (16, 28, 29) {real, imag} */,
  {32'hc36011db, 32'hc2e387d4} /* (16, 28, 28) {real, imag} */,
  {32'h42ce9854, 32'hc12498d6} /* (16, 28, 27) {real, imag} */,
  {32'h42f34626, 32'h424f4eb4} /* (16, 28, 26) {real, imag} */,
  {32'h42005a94, 32'hc27e4d84} /* (16, 28, 25) {real, imag} */,
  {32'hc223fe5e, 32'h42ad4b03} /* (16, 28, 24) {real, imag} */,
  {32'h4345c7e6, 32'h42658d25} /* (16, 28, 23) {real, imag} */,
  {32'hc21b2790, 32'hc1926d16} /* (16, 28, 22) {real, imag} */,
  {32'hc1c18860, 32'h4161b498} /* (16, 28, 21) {real, imag} */,
  {32'h41efa3ce, 32'hc3197897} /* (16, 28, 20) {real, imag} */,
  {32'h4246a6da, 32'hc06f6ee4} /* (16, 28, 19) {real, imag} */,
  {32'h41ed0e2c, 32'hc298b0d6} /* (16, 28, 18) {real, imag} */,
  {32'h3ef1b518, 32'h4228f16a} /* (16, 28, 17) {real, imag} */,
  {32'h4305d9d8, 32'h00000000} /* (16, 28, 16) {real, imag} */,
  {32'h3ef1b518, 32'hc228f16a} /* (16, 28, 15) {real, imag} */,
  {32'h41ed0e2c, 32'h4298b0d6} /* (16, 28, 14) {real, imag} */,
  {32'h4246a6da, 32'h406f6ee4} /* (16, 28, 13) {real, imag} */,
  {32'h41efa3ce, 32'h43197897} /* (16, 28, 12) {real, imag} */,
  {32'hc1c18860, 32'hc161b498} /* (16, 28, 11) {real, imag} */,
  {32'hc21b2790, 32'h41926d16} /* (16, 28, 10) {real, imag} */,
  {32'h4345c7e6, 32'hc2658d25} /* (16, 28, 9) {real, imag} */,
  {32'hc223fe5e, 32'hc2ad4b03} /* (16, 28, 8) {real, imag} */,
  {32'h42005a94, 32'h427e4d84} /* (16, 28, 7) {real, imag} */,
  {32'h42f34626, 32'hc24f4eb4} /* (16, 28, 6) {real, imag} */,
  {32'h42ce9854, 32'h412498d6} /* (16, 28, 5) {real, imag} */,
  {32'hc36011db, 32'h42e387d4} /* (16, 28, 4) {real, imag} */,
  {32'hc00235c8, 32'h4195f5be} /* (16, 28, 3) {real, imag} */,
  {32'h43dc085d, 32'h439cced3} /* (16, 28, 2) {real, imag} */,
  {32'hc4ca6a6d, 32'hc335b078} /* (16, 28, 1) {real, imag} */,
  {32'hc488915a, 32'h00000000} /* (16, 28, 0) {real, imag} */,
  {32'hc4b1f2a3, 32'h426199f0} /* (16, 27, 31) {real, imag} */,
  {32'h43b9beb0, 32'hc3570365} /* (16, 27, 30) {real, imag} */,
  {32'h4211121b, 32'hc107c53c} /* (16, 27, 29) {real, imag} */,
  {32'hc353ff3d, 32'hc28ad592} /* (16, 27, 28) {real, imag} */,
  {32'h42ded714, 32'h418efedc} /* (16, 27, 27) {real, imag} */,
  {32'h4298a654, 32'hc2b70b71} /* (16, 27, 26) {real, imag} */,
  {32'hc221cf64, 32'h41fd346c} /* (16, 27, 25) {real, imag} */,
  {32'hc2416f04, 32'hc22a26a6} /* (16, 27, 24) {real, imag} */,
  {32'h41c02bfd, 32'h4289c4d4} /* (16, 27, 23) {real, imag} */,
  {32'hc218a514, 32'hc2573e68} /* (16, 27, 22) {real, imag} */,
  {32'h40e38418, 32'hc24cf186} /* (16, 27, 21) {real, imag} */,
  {32'hc105916f, 32'hc234ceb7} /* (16, 27, 20) {real, imag} */,
  {32'h41a73c94, 32'h4289e064} /* (16, 27, 19) {real, imag} */,
  {32'h404ea2cc, 32'hbf3b5bb0} /* (16, 27, 18) {real, imag} */,
  {32'hc04d5ea8, 32'hc235d424} /* (16, 27, 17) {real, imag} */,
  {32'hc1853e48, 32'h00000000} /* (16, 27, 16) {real, imag} */,
  {32'hc04d5ea8, 32'h4235d424} /* (16, 27, 15) {real, imag} */,
  {32'h404ea2cc, 32'h3f3b5bb0} /* (16, 27, 14) {real, imag} */,
  {32'h41a73c94, 32'hc289e064} /* (16, 27, 13) {real, imag} */,
  {32'hc105916f, 32'h4234ceb7} /* (16, 27, 12) {real, imag} */,
  {32'h40e38418, 32'h424cf186} /* (16, 27, 11) {real, imag} */,
  {32'hc218a514, 32'h42573e68} /* (16, 27, 10) {real, imag} */,
  {32'h41c02bfd, 32'hc289c4d4} /* (16, 27, 9) {real, imag} */,
  {32'hc2416f04, 32'h422a26a6} /* (16, 27, 8) {real, imag} */,
  {32'hc221cf64, 32'hc1fd346c} /* (16, 27, 7) {real, imag} */,
  {32'h4298a654, 32'h42b70b71} /* (16, 27, 6) {real, imag} */,
  {32'h42ded714, 32'hc18efedc} /* (16, 27, 5) {real, imag} */,
  {32'hc353ff3d, 32'h428ad592} /* (16, 27, 4) {real, imag} */,
  {32'h4211121b, 32'h4107c53c} /* (16, 27, 3) {real, imag} */,
  {32'h43b9beb0, 32'h43570365} /* (16, 27, 2) {real, imag} */,
  {32'hc4b1f2a3, 32'hc26199f0} /* (16, 27, 1) {real, imag} */,
  {32'hc48cee4c, 32'h00000000} /* (16, 27, 0) {real, imag} */,
  {32'hc4a184df, 32'h3f16a200} /* (16, 26, 31) {real, imag} */,
  {32'h439e38cf, 32'hc30b80a2} /* (16, 26, 30) {real, imag} */,
  {32'h421a8528, 32'hc2567f06} /* (16, 26, 29) {real, imag} */,
  {32'hc36166a5, 32'hc2824484} /* (16, 26, 28) {real, imag} */,
  {32'h4182896a, 32'hc27aa0a8} /* (16, 26, 27) {real, imag} */,
  {32'h4275cd98, 32'hc27051e1} /* (16, 26, 26) {real, imag} */,
  {32'hc1bba58f, 32'hc1eb322f} /* (16, 26, 25) {real, imag} */,
  {32'h42512c32, 32'hc08ee860} /* (16, 26, 24) {real, imag} */,
  {32'h429e499f, 32'h408ffd6e} /* (16, 26, 23) {real, imag} */,
  {32'h42b48160, 32'h4258de66} /* (16, 26, 22) {real, imag} */,
  {32'h426ebc1c, 32'hc2e6bed2} /* (16, 26, 21) {real, imag} */,
  {32'hc28232fe, 32'hc12135c6} /* (16, 26, 20) {real, imag} */,
  {32'h41f61c06, 32'h423e6844} /* (16, 26, 19) {real, imag} */,
  {32'hc2296d25, 32'h418d8b4c} /* (16, 26, 18) {real, imag} */,
  {32'hc260f90f, 32'hc13cc277} /* (16, 26, 17) {real, imag} */,
  {32'hc1c2e71e, 32'h00000000} /* (16, 26, 16) {real, imag} */,
  {32'hc260f90f, 32'h413cc277} /* (16, 26, 15) {real, imag} */,
  {32'hc2296d25, 32'hc18d8b4c} /* (16, 26, 14) {real, imag} */,
  {32'h41f61c06, 32'hc23e6844} /* (16, 26, 13) {real, imag} */,
  {32'hc28232fe, 32'h412135c6} /* (16, 26, 12) {real, imag} */,
  {32'h426ebc1c, 32'h42e6bed2} /* (16, 26, 11) {real, imag} */,
  {32'h42b48160, 32'hc258de66} /* (16, 26, 10) {real, imag} */,
  {32'h429e499f, 32'hc08ffd6e} /* (16, 26, 9) {real, imag} */,
  {32'h42512c32, 32'h408ee860} /* (16, 26, 8) {real, imag} */,
  {32'hc1bba58f, 32'h41eb322f} /* (16, 26, 7) {real, imag} */,
  {32'h4275cd98, 32'h427051e1} /* (16, 26, 6) {real, imag} */,
  {32'h4182896a, 32'h427aa0a8} /* (16, 26, 5) {real, imag} */,
  {32'hc36166a5, 32'h42824484} /* (16, 26, 4) {real, imag} */,
  {32'h421a8528, 32'h42567f06} /* (16, 26, 3) {real, imag} */,
  {32'h439e38cf, 32'h430b80a2} /* (16, 26, 2) {real, imag} */,
  {32'hc4a184df, 32'hbf16a200} /* (16, 26, 1) {real, imag} */,
  {32'hc49e1ac1, 32'h00000000} /* (16, 26, 0) {real, imag} */,
  {32'hc49c833d, 32'h4292b61c} /* (16, 25, 31) {real, imag} */,
  {32'h439d580b, 32'hc302f988} /* (16, 25, 30) {real, imag} */,
  {32'hc1b4b334, 32'hc2d95ed9} /* (16, 25, 29) {real, imag} */,
  {32'hc345402c, 32'hc27d50e8} /* (16, 25, 28) {real, imag} */,
  {32'h432ae79d, 32'hc070c0c0} /* (16, 25, 27) {real, imag} */,
  {32'h4281f97c, 32'hc20eee40} /* (16, 25, 26) {real, imag} */,
  {32'hc2807510, 32'h3fd4ba70} /* (16, 25, 25) {real, imag} */,
  {32'h42d67009, 32'hc2944dd1} /* (16, 25, 24) {real, imag} */,
  {32'hc03cda20, 32'hc1f38b22} /* (16, 25, 23) {real, imag} */,
  {32'hc14a2f87, 32'h41d16af4} /* (16, 25, 22) {real, imag} */,
  {32'hc229f6a9, 32'hc23a6548} /* (16, 25, 21) {real, imag} */,
  {32'h422d6068, 32'hc290f5bd} /* (16, 25, 20) {real, imag} */,
  {32'h4250a6cc, 32'h42413074} /* (16, 25, 19) {real, imag} */,
  {32'hc17cad2c, 32'hc2253eaa} /* (16, 25, 18) {real, imag} */,
  {32'h42a8b1a0, 32'h42066b34} /* (16, 25, 17) {real, imag} */,
  {32'hc1eae242, 32'h00000000} /* (16, 25, 16) {real, imag} */,
  {32'h42a8b1a0, 32'hc2066b34} /* (16, 25, 15) {real, imag} */,
  {32'hc17cad2c, 32'h42253eaa} /* (16, 25, 14) {real, imag} */,
  {32'h4250a6cc, 32'hc2413074} /* (16, 25, 13) {real, imag} */,
  {32'h422d6068, 32'h4290f5bd} /* (16, 25, 12) {real, imag} */,
  {32'hc229f6a9, 32'h423a6548} /* (16, 25, 11) {real, imag} */,
  {32'hc14a2f87, 32'hc1d16af4} /* (16, 25, 10) {real, imag} */,
  {32'hc03cda20, 32'h41f38b22} /* (16, 25, 9) {real, imag} */,
  {32'h42d67009, 32'h42944dd1} /* (16, 25, 8) {real, imag} */,
  {32'hc2807510, 32'hbfd4ba70} /* (16, 25, 7) {real, imag} */,
  {32'h4281f97c, 32'h420eee40} /* (16, 25, 6) {real, imag} */,
  {32'h432ae79d, 32'h4070c0c0} /* (16, 25, 5) {real, imag} */,
  {32'hc345402c, 32'h427d50e8} /* (16, 25, 4) {real, imag} */,
  {32'hc1b4b334, 32'h42d95ed9} /* (16, 25, 3) {real, imag} */,
  {32'h439d580b, 32'h4302f988} /* (16, 25, 2) {real, imag} */,
  {32'hc49c833d, 32'hc292b61c} /* (16, 25, 1) {real, imag} */,
  {32'hc49956ac, 32'h00000000} /* (16, 25, 0) {real, imag} */,
  {32'hc48e3966, 32'h42a58e50} /* (16, 24, 31) {real, imag} */,
  {32'h43df03d2, 32'hc34f4914} /* (16, 24, 30) {real, imag} */,
  {32'hc24e02dc, 32'hc336c37d} /* (16, 24, 29) {real, imag} */,
  {32'hc383d40f, 32'hc2bc08b0} /* (16, 24, 28) {real, imag} */,
  {32'h431fbac6, 32'hc2ff6ca8} /* (16, 24, 27) {real, imag} */,
  {32'h426cef47, 32'h42960c67} /* (16, 24, 26) {real, imag} */,
  {32'hc2bf16ce, 32'hc1d32bba} /* (16, 24, 25) {real, imag} */,
  {32'h42e2485e, 32'hc1676554} /* (16, 24, 24) {real, imag} */,
  {32'h42cce6e3, 32'h429c21fb} /* (16, 24, 23) {real, imag} */,
  {32'h425d3fe1, 32'h4211291c} /* (16, 24, 22) {real, imag} */,
  {32'h41915964, 32'hc1f29743} /* (16, 24, 21) {real, imag} */,
  {32'h41714dc0, 32'h42a63bca} /* (16, 24, 20) {real, imag} */,
  {32'hc242ffc1, 32'hc206adae} /* (16, 24, 19) {real, imag} */,
  {32'h422d1f3e, 32'h42948f54} /* (16, 24, 18) {real, imag} */,
  {32'h420ac37e, 32'hc2a7912a} /* (16, 24, 17) {real, imag} */,
  {32'h4255196c, 32'h00000000} /* (16, 24, 16) {real, imag} */,
  {32'h420ac37e, 32'h42a7912a} /* (16, 24, 15) {real, imag} */,
  {32'h422d1f3e, 32'hc2948f54} /* (16, 24, 14) {real, imag} */,
  {32'hc242ffc1, 32'h4206adae} /* (16, 24, 13) {real, imag} */,
  {32'h41714dc0, 32'hc2a63bca} /* (16, 24, 12) {real, imag} */,
  {32'h41915964, 32'h41f29743} /* (16, 24, 11) {real, imag} */,
  {32'h425d3fe1, 32'hc211291c} /* (16, 24, 10) {real, imag} */,
  {32'h42cce6e3, 32'hc29c21fb} /* (16, 24, 9) {real, imag} */,
  {32'h42e2485e, 32'h41676554} /* (16, 24, 8) {real, imag} */,
  {32'hc2bf16ce, 32'h41d32bba} /* (16, 24, 7) {real, imag} */,
  {32'h426cef47, 32'hc2960c67} /* (16, 24, 6) {real, imag} */,
  {32'h431fbac6, 32'h42ff6ca8} /* (16, 24, 5) {real, imag} */,
  {32'hc383d40f, 32'h42bc08b0} /* (16, 24, 4) {real, imag} */,
  {32'hc24e02dc, 32'h4336c37d} /* (16, 24, 3) {real, imag} */,
  {32'h43df03d2, 32'h434f4914} /* (16, 24, 2) {real, imag} */,
  {32'hc48e3966, 32'hc2a58e50} /* (16, 24, 1) {real, imag} */,
  {32'hc497702b, 32'h00000000} /* (16, 24, 0) {real, imag} */,
  {32'hc4565dea, 32'h4301d4de} /* (16, 23, 31) {real, imag} */,
  {32'h43fbefd7, 32'hc1d31a21} /* (16, 23, 30) {real, imag} */,
  {32'hc275cf7b, 32'hc2e7c415} /* (16, 23, 29) {real, imag} */,
  {32'hc3469827, 32'hc300f6b7} /* (16, 23, 28) {real, imag} */,
  {32'h429599b2, 32'hc26bd2d8} /* (16, 23, 27) {real, imag} */,
  {32'hc303639f, 32'hc24a62dc} /* (16, 23, 26) {real, imag} */,
  {32'hc30b5e03, 32'h40bb09a8} /* (16, 23, 25) {real, imag} */,
  {32'h4316476d, 32'hc245650e} /* (16, 23, 24) {real, imag} */,
  {32'h42d2b543, 32'hc214449d} /* (16, 23, 23) {real, imag} */,
  {32'h42aa3cbb, 32'hc23eaffe} /* (16, 23, 22) {real, imag} */,
  {32'h422e4734, 32'h42ae8eb7} /* (16, 23, 21) {real, imag} */,
  {32'hc29474c2, 32'h42bb0cc4} /* (16, 23, 20) {real, imag} */,
  {32'h41e8ebec, 32'h4061d080} /* (16, 23, 19) {real, imag} */,
  {32'hbebdd700, 32'hc2e62c15} /* (16, 23, 18) {real, imag} */,
  {32'hc22bcd02, 32'h4237dadd} /* (16, 23, 17) {real, imag} */,
  {32'h425c2aaa, 32'h00000000} /* (16, 23, 16) {real, imag} */,
  {32'hc22bcd02, 32'hc237dadd} /* (16, 23, 15) {real, imag} */,
  {32'hbebdd700, 32'h42e62c15} /* (16, 23, 14) {real, imag} */,
  {32'h41e8ebec, 32'hc061d080} /* (16, 23, 13) {real, imag} */,
  {32'hc29474c2, 32'hc2bb0cc4} /* (16, 23, 12) {real, imag} */,
  {32'h422e4734, 32'hc2ae8eb7} /* (16, 23, 11) {real, imag} */,
  {32'h42aa3cbb, 32'h423eaffe} /* (16, 23, 10) {real, imag} */,
  {32'h42d2b543, 32'h4214449d} /* (16, 23, 9) {real, imag} */,
  {32'h4316476d, 32'h4245650e} /* (16, 23, 8) {real, imag} */,
  {32'hc30b5e03, 32'hc0bb09a8} /* (16, 23, 7) {real, imag} */,
  {32'hc303639f, 32'h424a62dc} /* (16, 23, 6) {real, imag} */,
  {32'h429599b2, 32'h426bd2d8} /* (16, 23, 5) {real, imag} */,
  {32'hc3469827, 32'h4300f6b7} /* (16, 23, 4) {real, imag} */,
  {32'hc275cf7b, 32'h42e7c415} /* (16, 23, 3) {real, imag} */,
  {32'h43fbefd7, 32'h41d31a21} /* (16, 23, 2) {real, imag} */,
  {32'hc4565dea, 32'hc301d4de} /* (16, 23, 1) {real, imag} */,
  {32'hc489fc32, 32'h00000000} /* (16, 23, 0) {real, imag} */,
  {32'hc4372cca, 32'h42b95010} /* (16, 22, 31) {real, imag} */,
  {32'h43cb5dfa, 32'hc1c92c7a} /* (16, 22, 30) {real, imag} */,
  {32'hc2846ed6, 32'hc23adec2} /* (16, 22, 29) {real, imag} */,
  {32'hc33ec336, 32'hc27e2b93} /* (16, 22, 28) {real, imag} */,
  {32'h42aedfa6, 32'hc1dda36d} /* (16, 22, 27) {real, imag} */,
  {32'hc0ed23c8, 32'hc2906468} /* (16, 22, 26) {real, imag} */,
  {32'h419f90e5, 32'h427e6dbe} /* (16, 22, 25) {real, imag} */,
  {32'h42135044, 32'hc1f723cc} /* (16, 22, 24) {real, imag} */,
  {32'hc23f3062, 32'hc26d3314} /* (16, 22, 23) {real, imag} */,
  {32'h4210b2f2, 32'h42a71cae} /* (16, 22, 22) {real, imag} */,
  {32'hc174f177, 32'hc29bcfcc} /* (16, 22, 21) {real, imag} */,
  {32'h427d2c05, 32'hc21e6a70} /* (16, 22, 20) {real, imag} */,
  {32'h425c6dae, 32'h421f680a} /* (16, 22, 19) {real, imag} */,
  {32'h42802e00, 32'hc242e1d1} /* (16, 22, 18) {real, imag} */,
  {32'h42463f2c, 32'h425a0fb4} /* (16, 22, 17) {real, imag} */,
  {32'h4106acd8, 32'h00000000} /* (16, 22, 16) {real, imag} */,
  {32'h42463f2c, 32'hc25a0fb4} /* (16, 22, 15) {real, imag} */,
  {32'h42802e00, 32'h4242e1d1} /* (16, 22, 14) {real, imag} */,
  {32'h425c6dae, 32'hc21f680a} /* (16, 22, 13) {real, imag} */,
  {32'h427d2c05, 32'h421e6a70} /* (16, 22, 12) {real, imag} */,
  {32'hc174f177, 32'h429bcfcc} /* (16, 22, 11) {real, imag} */,
  {32'h4210b2f2, 32'hc2a71cae} /* (16, 22, 10) {real, imag} */,
  {32'hc23f3062, 32'h426d3314} /* (16, 22, 9) {real, imag} */,
  {32'h42135044, 32'h41f723cc} /* (16, 22, 8) {real, imag} */,
  {32'h419f90e5, 32'hc27e6dbe} /* (16, 22, 7) {real, imag} */,
  {32'hc0ed23c8, 32'h42906468} /* (16, 22, 6) {real, imag} */,
  {32'h42aedfa6, 32'h41dda36d} /* (16, 22, 5) {real, imag} */,
  {32'hc33ec336, 32'h427e2b93} /* (16, 22, 4) {real, imag} */,
  {32'hc2846ed6, 32'h423adec2} /* (16, 22, 3) {real, imag} */,
  {32'h43cb5dfa, 32'h41c92c7a} /* (16, 22, 2) {real, imag} */,
  {32'hc4372cca, 32'hc2b95010} /* (16, 22, 1) {real, imag} */,
  {32'hc46f4ab9, 32'h00000000} /* (16, 22, 0) {real, imag} */,
  {32'hc3a7658a, 32'h423eace0} /* (16, 21, 31) {real, imag} */,
  {32'h437ddfe0, 32'h42a8de70} /* (16, 21, 30) {real, imag} */,
  {32'h4282a200, 32'hc0ea8168} /* (16, 21, 29) {real, imag} */,
  {32'h4230c732, 32'hc2b4c189} /* (16, 21, 28) {real, imag} */,
  {32'hc1cb4ed0, 32'hc1aceee1} /* (16, 21, 27) {real, imag} */,
  {32'h41b1c8c6, 32'hc2209e7c} /* (16, 21, 26) {real, imag} */,
  {32'h42bf34c8, 32'h42826530} /* (16, 21, 25) {real, imag} */,
  {32'hc09deefc, 32'hc285c282} /* (16, 21, 24) {real, imag} */,
  {32'h41990fd1, 32'h42800618} /* (16, 21, 23) {real, imag} */,
  {32'h410954c0, 32'h428e46c0} /* (16, 21, 22) {real, imag} */,
  {32'hc2afcdac, 32'h420479f0} /* (16, 21, 21) {real, imag} */,
  {32'hc2bbd1e8, 32'h3fed7ae0} /* (16, 21, 20) {real, imag} */,
  {32'hbfada2e0, 32'hc2930e2d} /* (16, 21, 19) {real, imag} */,
  {32'h418d04b4, 32'h42248835} /* (16, 21, 18) {real, imag} */,
  {32'h41fd1873, 32'hc2677525} /* (16, 21, 17) {real, imag} */,
  {32'hc06ef940, 32'h00000000} /* (16, 21, 16) {real, imag} */,
  {32'h41fd1873, 32'h42677525} /* (16, 21, 15) {real, imag} */,
  {32'h418d04b4, 32'hc2248835} /* (16, 21, 14) {real, imag} */,
  {32'hbfada2e0, 32'h42930e2d} /* (16, 21, 13) {real, imag} */,
  {32'hc2bbd1e8, 32'hbfed7ae0} /* (16, 21, 12) {real, imag} */,
  {32'hc2afcdac, 32'hc20479f0} /* (16, 21, 11) {real, imag} */,
  {32'h410954c0, 32'hc28e46c0} /* (16, 21, 10) {real, imag} */,
  {32'h41990fd1, 32'hc2800618} /* (16, 21, 9) {real, imag} */,
  {32'hc09deefc, 32'h4285c282} /* (16, 21, 8) {real, imag} */,
  {32'h42bf34c8, 32'hc2826530} /* (16, 21, 7) {real, imag} */,
  {32'h41b1c8c6, 32'h42209e7c} /* (16, 21, 6) {real, imag} */,
  {32'hc1cb4ed0, 32'h41aceee1} /* (16, 21, 5) {real, imag} */,
  {32'h4230c732, 32'h42b4c189} /* (16, 21, 4) {real, imag} */,
  {32'h4282a200, 32'h40ea8168} /* (16, 21, 3) {real, imag} */,
  {32'h437ddfe0, 32'hc2a8de70} /* (16, 21, 2) {real, imag} */,
  {32'hc3a7658a, 32'hc23eace0} /* (16, 21, 1) {real, imag} */,
  {32'hc42bf9d9, 32'h00000000} /* (16, 21, 0) {real, imag} */,
  {32'h438408a5, 32'h42148354} /* (16, 20, 31) {real, imag} */,
  {32'hc152aeb0, 32'h435b1b6e} /* (16, 20, 30) {real, imag} */,
  {32'h420fc4dc, 32'h42de8461} /* (16, 20, 29) {real, imag} */,
  {32'h435a4586, 32'hc2f9181f} /* (16, 20, 28) {real, imag} */,
  {32'hc2e39916, 32'h4132ba48} /* (16, 20, 27) {real, imag} */,
  {32'hc3538d6c, 32'hc30152f2} /* (16, 20, 26) {real, imag} */,
  {32'h422b4658, 32'h41bc11d2} /* (16, 20, 25) {real, imag} */,
  {32'hc2e3e9a6, 32'h403190e0} /* (16, 20, 24) {real, imag} */,
  {32'h414ec188, 32'hc1368010} /* (16, 20, 23) {real, imag} */,
  {32'hc2a6af60, 32'hc214e9e8} /* (16, 20, 22) {real, imag} */,
  {32'h42b50792, 32'hc1d15554} /* (16, 20, 21) {real, imag} */,
  {32'h420f4888, 32'h40cb62c8} /* (16, 20, 20) {real, imag} */,
  {32'hc21337b2, 32'hc0645ef8} /* (16, 20, 19) {real, imag} */,
  {32'h41d1117e, 32'hc09b49c0} /* (16, 20, 18) {real, imag} */,
  {32'h4283ba0a, 32'h42448a7c} /* (16, 20, 17) {real, imag} */,
  {32'h40f02ccc, 32'h00000000} /* (16, 20, 16) {real, imag} */,
  {32'h4283ba0a, 32'hc2448a7c} /* (16, 20, 15) {real, imag} */,
  {32'h41d1117e, 32'h409b49c0} /* (16, 20, 14) {real, imag} */,
  {32'hc21337b2, 32'h40645ef8} /* (16, 20, 13) {real, imag} */,
  {32'h420f4888, 32'hc0cb62c8} /* (16, 20, 12) {real, imag} */,
  {32'h42b50792, 32'h41d15554} /* (16, 20, 11) {real, imag} */,
  {32'hc2a6af60, 32'h4214e9e8} /* (16, 20, 10) {real, imag} */,
  {32'h414ec188, 32'h41368010} /* (16, 20, 9) {real, imag} */,
  {32'hc2e3e9a6, 32'hc03190e0} /* (16, 20, 8) {real, imag} */,
  {32'h422b4658, 32'hc1bc11d2} /* (16, 20, 7) {real, imag} */,
  {32'hc3538d6c, 32'h430152f2} /* (16, 20, 6) {real, imag} */,
  {32'hc2e39916, 32'hc132ba48} /* (16, 20, 5) {real, imag} */,
  {32'h435a4586, 32'h42f9181f} /* (16, 20, 4) {real, imag} */,
  {32'h420fc4dc, 32'hc2de8461} /* (16, 20, 3) {real, imag} */,
  {32'hc152aeb0, 32'hc35b1b6e} /* (16, 20, 2) {real, imag} */,
  {32'h438408a5, 32'hc2148354} /* (16, 20, 1) {real, imag} */,
  {32'hc10fc120, 32'h00000000} /* (16, 20, 0) {real, imag} */,
  {32'h440582e0, 32'h3fbb1700} /* (16, 19, 31) {real, imag} */,
  {32'hc366c1d1, 32'h438d33e5} /* (16, 19, 30) {real, imag} */,
  {32'h4342ebed, 32'h42c8f931} /* (16, 19, 29) {real, imag} */,
  {32'h43178a0c, 32'hc17fde90} /* (16, 19, 28) {real, imag} */,
  {32'hc32fb97e, 32'h42237cdc} /* (16, 19, 27) {real, imag} */,
  {32'h422b9a48, 32'h42a321b2} /* (16, 19, 26) {real, imag} */,
  {32'h4305ccab, 32'hc2b80055} /* (16, 19, 25) {real, imag} */,
  {32'hc2e112fc, 32'h432da6b8} /* (16, 19, 24) {real, imag} */,
  {32'hc0bec778, 32'h41df7e08} /* (16, 19, 23) {real, imag} */,
  {32'hc0da0af0, 32'hc1055543} /* (16, 19, 22) {real, imag} */,
  {32'h41a71f6c, 32'h41cbd870} /* (16, 19, 21) {real, imag} */,
  {32'hc2c2cb54, 32'hc0460230} /* (16, 19, 20) {real, imag} */,
  {32'h421abdb1, 32'h40b12781} /* (16, 19, 19) {real, imag} */,
  {32'hc20b3b3c, 32'h420a2f9e} /* (16, 19, 18) {real, imag} */,
  {32'hc21b0cb2, 32'h41eae296} /* (16, 19, 17) {real, imag} */,
  {32'h41e549e4, 32'h00000000} /* (16, 19, 16) {real, imag} */,
  {32'hc21b0cb2, 32'hc1eae296} /* (16, 19, 15) {real, imag} */,
  {32'hc20b3b3c, 32'hc20a2f9e} /* (16, 19, 14) {real, imag} */,
  {32'h421abdb1, 32'hc0b12781} /* (16, 19, 13) {real, imag} */,
  {32'hc2c2cb54, 32'h40460230} /* (16, 19, 12) {real, imag} */,
  {32'h41a71f6c, 32'hc1cbd870} /* (16, 19, 11) {real, imag} */,
  {32'hc0da0af0, 32'h41055543} /* (16, 19, 10) {real, imag} */,
  {32'hc0bec778, 32'hc1df7e08} /* (16, 19, 9) {real, imag} */,
  {32'hc2e112fc, 32'hc32da6b8} /* (16, 19, 8) {real, imag} */,
  {32'h4305ccab, 32'h42b80055} /* (16, 19, 7) {real, imag} */,
  {32'h422b9a48, 32'hc2a321b2} /* (16, 19, 6) {real, imag} */,
  {32'hc32fb97e, 32'hc2237cdc} /* (16, 19, 5) {real, imag} */,
  {32'h43178a0c, 32'h417fde90} /* (16, 19, 4) {real, imag} */,
  {32'h4342ebed, 32'hc2c8f931} /* (16, 19, 3) {real, imag} */,
  {32'hc366c1d1, 32'hc38d33e5} /* (16, 19, 2) {real, imag} */,
  {32'h440582e0, 32'hbfbb1700} /* (16, 19, 1) {real, imag} */,
  {32'h43c3540e, 32'h00000000} /* (16, 19, 0) {real, imag} */,
  {32'h444aa1e0, 32'hc2887656} /* (16, 18, 31) {real, imag} */,
  {32'hc3efc907, 32'h42ac0464} /* (16, 18, 30) {real, imag} */,
  {32'h4382d715, 32'h430cf94c} /* (16, 18, 29) {real, imag} */,
  {32'h43183d4a, 32'h41e336e8} /* (16, 18, 28) {real, imag} */,
  {32'hc279c3bc, 32'h423e6b74} /* (16, 18, 27) {real, imag} */,
  {32'h421598ac, 32'hc2903a11} /* (16, 18, 26) {real, imag} */,
  {32'h42c2ac2a, 32'h42266f57} /* (16, 18, 25) {real, imag} */,
  {32'h41a06d8a, 32'hc19e2e14} /* (16, 18, 24) {real, imag} */,
  {32'hc2b3fb90, 32'h414c8b3e} /* (16, 18, 23) {real, imag} */,
  {32'hc24893b9, 32'h42c23642} /* (16, 18, 22) {real, imag} */,
  {32'h42308db5, 32'h42cf92da} /* (16, 18, 21) {real, imag} */,
  {32'hc245496e, 32'hc1c7a834} /* (16, 18, 20) {real, imag} */,
  {32'hc2d229dc, 32'hc2a3f59a} /* (16, 18, 19) {real, imag} */,
  {32'h40fc7e4e, 32'h425563e0} /* (16, 18, 18) {real, imag} */,
  {32'hc1995f8e, 32'hc21d4840} /* (16, 18, 17) {real, imag} */,
  {32'h425c474c, 32'h00000000} /* (16, 18, 16) {real, imag} */,
  {32'hc1995f8e, 32'h421d4840} /* (16, 18, 15) {real, imag} */,
  {32'h40fc7e4e, 32'hc25563e0} /* (16, 18, 14) {real, imag} */,
  {32'hc2d229dc, 32'h42a3f59a} /* (16, 18, 13) {real, imag} */,
  {32'hc245496e, 32'h41c7a834} /* (16, 18, 12) {real, imag} */,
  {32'h42308db5, 32'hc2cf92da} /* (16, 18, 11) {real, imag} */,
  {32'hc24893b9, 32'hc2c23642} /* (16, 18, 10) {real, imag} */,
  {32'hc2b3fb90, 32'hc14c8b3e} /* (16, 18, 9) {real, imag} */,
  {32'h41a06d8a, 32'h419e2e14} /* (16, 18, 8) {real, imag} */,
  {32'h42c2ac2a, 32'hc2266f57} /* (16, 18, 7) {real, imag} */,
  {32'h421598ac, 32'h42903a11} /* (16, 18, 6) {real, imag} */,
  {32'hc279c3bc, 32'hc23e6b74} /* (16, 18, 5) {real, imag} */,
  {32'h43183d4a, 32'hc1e336e8} /* (16, 18, 4) {real, imag} */,
  {32'h4382d715, 32'hc30cf94c} /* (16, 18, 3) {real, imag} */,
  {32'hc3efc907, 32'hc2ac0464} /* (16, 18, 2) {real, imag} */,
  {32'h444aa1e0, 32'h42887656} /* (16, 18, 1) {real, imag} */,
  {32'h442d92d1, 32'h00000000} /* (16, 18, 0) {real, imag} */,
  {32'h446a1dd3, 32'hc2e1133c} /* (16, 17, 31) {real, imag} */,
  {32'hc4197ade, 32'h427af27a} /* (16, 17, 30) {real, imag} */,
  {32'h439262bc, 32'hc2a2c4d9} /* (16, 17, 29) {real, imag} */,
  {32'h433addec, 32'h42a2e3b7} /* (16, 17, 28) {real, imag} */,
  {32'hc302bc64, 32'h415eeac8} /* (16, 17, 27) {real, imag} */,
  {32'hc0c1fde0, 32'hc2e68f96} /* (16, 17, 26) {real, imag} */,
  {32'h422a47e5, 32'hc2b2e06d} /* (16, 17, 25) {real, imag} */,
  {32'h42e86a29, 32'h42ae4683} /* (16, 17, 24) {real, imag} */,
  {32'h42ba7213, 32'hc1b2f2e0} /* (16, 17, 23) {real, imag} */,
  {32'hbfb855d0, 32'hc3055af8} /* (16, 17, 22) {real, imag} */,
  {32'hc28d89fe, 32'h4322673e} /* (16, 17, 21) {real, imag} */,
  {32'h4233a17f, 32'h4298e397} /* (16, 17, 20) {real, imag} */,
  {32'hc2305122, 32'hc23c2f19} /* (16, 17, 19) {real, imag} */,
  {32'hc220a2f6, 32'h42462c5d} /* (16, 17, 18) {real, imag} */,
  {32'h41fb4642, 32'h3ed600c0} /* (16, 17, 17) {real, imag} */,
  {32'h41f80378, 32'h00000000} /* (16, 17, 16) {real, imag} */,
  {32'h41fb4642, 32'hbed600c0} /* (16, 17, 15) {real, imag} */,
  {32'hc220a2f6, 32'hc2462c5d} /* (16, 17, 14) {real, imag} */,
  {32'hc2305122, 32'h423c2f19} /* (16, 17, 13) {real, imag} */,
  {32'h4233a17f, 32'hc298e397} /* (16, 17, 12) {real, imag} */,
  {32'hc28d89fe, 32'hc322673e} /* (16, 17, 11) {real, imag} */,
  {32'hbfb855d0, 32'h43055af8} /* (16, 17, 10) {real, imag} */,
  {32'h42ba7213, 32'h41b2f2e0} /* (16, 17, 9) {real, imag} */,
  {32'h42e86a29, 32'hc2ae4683} /* (16, 17, 8) {real, imag} */,
  {32'h422a47e5, 32'h42b2e06d} /* (16, 17, 7) {real, imag} */,
  {32'hc0c1fde0, 32'h42e68f96} /* (16, 17, 6) {real, imag} */,
  {32'hc302bc64, 32'hc15eeac8} /* (16, 17, 5) {real, imag} */,
  {32'h433addec, 32'hc2a2e3b7} /* (16, 17, 4) {real, imag} */,
  {32'h439262bc, 32'h42a2c4d9} /* (16, 17, 3) {real, imag} */,
  {32'hc4197ade, 32'hc27af27a} /* (16, 17, 2) {real, imag} */,
  {32'h446a1dd3, 32'h42e1133c} /* (16, 17, 1) {real, imag} */,
  {32'h4436565e, 32'h00000000} /* (16, 17, 0) {real, imag} */,
  {32'h44780559, 32'hc20296a0} /* (16, 16, 31) {real, imag} */,
  {32'hc401073f, 32'h42ad03ca} /* (16, 16, 30) {real, imag} */,
  {32'h430b83d3, 32'hc28a6e34} /* (16, 16, 29) {real, imag} */,
  {32'h42ddeeb9, 32'h42a13f5b} /* (16, 16, 28) {real, imag} */,
  {32'hc35c9e1d, 32'h4321a39e} /* (16, 16, 27) {real, imag} */,
  {32'hc26a7d40, 32'h41a5ef96} /* (16, 16, 26) {real, imag} */,
  {32'h429b5a23, 32'hc1bba47e} /* (16, 16, 25) {real, imag} */,
  {32'hc0e42a40, 32'h4005a5c0} /* (16, 16, 24) {real, imag} */,
  {32'h41fcd110, 32'hc2277a71} /* (16, 16, 23) {real, imag} */,
  {32'hc1ceb671, 32'hc2173899} /* (16, 16, 22) {real, imag} */,
  {32'hc2bf7a77, 32'h41f03dc4} /* (16, 16, 21) {real, imag} */,
  {32'h4289d87e, 32'hc3164d26} /* (16, 16, 20) {real, imag} */,
  {32'h427318ae, 32'h423b1f50} /* (16, 16, 19) {real, imag} */,
  {32'hc2bff628, 32'hc203c9ea} /* (16, 16, 18) {real, imag} */,
  {32'h41855448, 32'h41a33db3} /* (16, 16, 17) {real, imag} */,
  {32'hc2221375, 32'h00000000} /* (16, 16, 16) {real, imag} */,
  {32'h41855448, 32'hc1a33db3} /* (16, 16, 15) {real, imag} */,
  {32'hc2bff628, 32'h4203c9ea} /* (16, 16, 14) {real, imag} */,
  {32'h427318ae, 32'hc23b1f50} /* (16, 16, 13) {real, imag} */,
  {32'h4289d87e, 32'h43164d26} /* (16, 16, 12) {real, imag} */,
  {32'hc2bf7a77, 32'hc1f03dc4} /* (16, 16, 11) {real, imag} */,
  {32'hc1ceb671, 32'h42173899} /* (16, 16, 10) {real, imag} */,
  {32'h41fcd110, 32'h42277a71} /* (16, 16, 9) {real, imag} */,
  {32'hc0e42a40, 32'hc005a5c0} /* (16, 16, 8) {real, imag} */,
  {32'h429b5a23, 32'h41bba47e} /* (16, 16, 7) {real, imag} */,
  {32'hc26a7d40, 32'hc1a5ef96} /* (16, 16, 6) {real, imag} */,
  {32'hc35c9e1d, 32'hc321a39e} /* (16, 16, 5) {real, imag} */,
  {32'h42ddeeb9, 32'hc2a13f5b} /* (16, 16, 4) {real, imag} */,
  {32'h430b83d3, 32'h428a6e34} /* (16, 16, 3) {real, imag} */,
  {32'hc401073f, 32'hc2ad03ca} /* (16, 16, 2) {real, imag} */,
  {32'h44780559, 32'h420296a0} /* (16, 16, 1) {real, imag} */,
  {32'h44047db0, 32'h00000000} /* (16, 16, 0) {real, imag} */,
  {32'h444df0f1, 32'h432cfd26} /* (16, 15, 31) {real, imag} */,
  {32'hc3e9459c, 32'h422955b6} /* (16, 15, 30) {real, imag} */,
  {32'h4317a0aa, 32'hc28a6d39} /* (16, 15, 29) {real, imag} */,
  {32'hc2467be6, 32'h43025c90} /* (16, 15, 28) {real, imag} */,
  {32'hc349b074, 32'h4307b424} /* (16, 15, 27) {real, imag} */,
  {32'h41b84f22, 32'h42aaf756} /* (16, 15, 26) {real, imag} */,
  {32'h4194f55a, 32'hc29d436b} /* (16, 15, 25) {real, imag} */,
  {32'hc1b2c324, 32'h410fef68} /* (16, 15, 24) {real, imag} */,
  {32'h419c2ebc, 32'h3eeab7a0} /* (16, 15, 23) {real, imag} */,
  {32'h426ef5aa, 32'hc22a047e} /* (16, 15, 22) {real, imag} */,
  {32'hc1e3e8df, 32'h420dceaa} /* (16, 15, 21) {real, imag} */,
  {32'hc2768e75, 32'h3fee1500} /* (16, 15, 20) {real, imag} */,
  {32'hc1865981, 32'hc148ca70} /* (16, 15, 19) {real, imag} */,
  {32'h41d96cc9, 32'hbffc7420} /* (16, 15, 18) {real, imag} */,
  {32'h4107ab4c, 32'h424d19a0} /* (16, 15, 17) {real, imag} */,
  {32'hc111c2f1, 32'h00000000} /* (16, 15, 16) {real, imag} */,
  {32'h4107ab4c, 32'hc24d19a0} /* (16, 15, 15) {real, imag} */,
  {32'h41d96cc9, 32'h3ffc7420} /* (16, 15, 14) {real, imag} */,
  {32'hc1865981, 32'h4148ca70} /* (16, 15, 13) {real, imag} */,
  {32'hc2768e75, 32'hbfee1500} /* (16, 15, 12) {real, imag} */,
  {32'hc1e3e8df, 32'hc20dceaa} /* (16, 15, 11) {real, imag} */,
  {32'h426ef5aa, 32'h422a047e} /* (16, 15, 10) {real, imag} */,
  {32'h419c2ebc, 32'hbeeab7a0} /* (16, 15, 9) {real, imag} */,
  {32'hc1b2c324, 32'hc10fef68} /* (16, 15, 8) {real, imag} */,
  {32'h4194f55a, 32'h429d436b} /* (16, 15, 7) {real, imag} */,
  {32'h41b84f22, 32'hc2aaf756} /* (16, 15, 6) {real, imag} */,
  {32'hc349b074, 32'hc307b424} /* (16, 15, 5) {real, imag} */,
  {32'hc2467be6, 32'hc3025c90} /* (16, 15, 4) {real, imag} */,
  {32'h4317a0aa, 32'h428a6d39} /* (16, 15, 3) {real, imag} */,
  {32'hc3e9459c, 32'hc22955b6} /* (16, 15, 2) {real, imag} */,
  {32'h444df0f1, 32'hc32cfd26} /* (16, 15, 1) {real, imag} */,
  {32'h4422978e, 32'h00000000} /* (16, 15, 0) {real, imag} */,
  {32'h4424a678, 32'h4339e65d} /* (16, 14, 31) {real, imag} */,
  {32'hc3bf37d1, 32'h42a64b56} /* (16, 14, 30) {real, imag} */,
  {32'h42a13704, 32'h41014ec0} /* (16, 14, 29) {real, imag} */,
  {32'h42a76594, 32'h41863b48} /* (16, 14, 28) {real, imag} */,
  {32'hc386629a, 32'h42134048} /* (16, 14, 27) {real, imag} */,
  {32'h42857a2a, 32'h41984c2f} /* (16, 14, 26) {real, imag} */,
  {32'h41cd4360, 32'hc30003e4} /* (16, 14, 25) {real, imag} */,
  {32'hc28f32ba, 32'h4236433a} /* (16, 14, 24) {real, imag} */,
  {32'h41c90014, 32'hc0980a7d} /* (16, 14, 23) {real, imag} */,
  {32'hc0a73728, 32'h415a7d30} /* (16, 14, 22) {real, imag} */,
  {32'h428a500a, 32'h4213d935} /* (16, 14, 21) {real, imag} */,
  {32'h4002c1e8, 32'hc01b72d0} /* (16, 14, 20) {real, imag} */,
  {32'h42445da4, 32'hc199e345} /* (16, 14, 19) {real, imag} */,
  {32'hc201e688, 32'hc1f6b6d0} /* (16, 14, 18) {real, imag} */,
  {32'hc273f7a3, 32'hc1af9af3} /* (16, 14, 17) {real, imag} */,
  {32'hc175fa00, 32'h00000000} /* (16, 14, 16) {real, imag} */,
  {32'hc273f7a3, 32'h41af9af3} /* (16, 14, 15) {real, imag} */,
  {32'hc201e688, 32'h41f6b6d0} /* (16, 14, 14) {real, imag} */,
  {32'h42445da4, 32'h4199e345} /* (16, 14, 13) {real, imag} */,
  {32'h4002c1e8, 32'h401b72d0} /* (16, 14, 12) {real, imag} */,
  {32'h428a500a, 32'hc213d935} /* (16, 14, 11) {real, imag} */,
  {32'hc0a73728, 32'hc15a7d30} /* (16, 14, 10) {real, imag} */,
  {32'h41c90014, 32'h40980a7d} /* (16, 14, 9) {real, imag} */,
  {32'hc28f32ba, 32'hc236433a} /* (16, 14, 8) {real, imag} */,
  {32'h41cd4360, 32'h430003e4} /* (16, 14, 7) {real, imag} */,
  {32'h42857a2a, 32'hc1984c2f} /* (16, 14, 6) {real, imag} */,
  {32'hc386629a, 32'hc2134048} /* (16, 14, 5) {real, imag} */,
  {32'h42a76594, 32'hc1863b48} /* (16, 14, 4) {real, imag} */,
  {32'h42a13704, 32'hc1014ec0} /* (16, 14, 3) {real, imag} */,
  {32'hc3bf37d1, 32'hc2a64b56} /* (16, 14, 2) {real, imag} */,
  {32'h4424a678, 32'hc339e65d} /* (16, 14, 1) {real, imag} */,
  {32'h4415a1cb, 32'h00000000} /* (16, 14, 0) {real, imag} */,
  {32'h442bb184, 32'h43455032} /* (16, 13, 31) {real, imag} */,
  {32'hc3a33508, 32'h42a01623} /* (16, 13, 30) {real, imag} */,
  {32'hc2537f90, 32'h42418122} /* (16, 13, 29) {real, imag} */,
  {32'h42e219a8, 32'h42c0a6aa} /* (16, 13, 28) {real, imag} */,
  {32'hc345b854, 32'h4200665c} /* (16, 13, 27) {real, imag} */,
  {32'hc2b31e6e, 32'hc1d655fa} /* (16, 13, 26) {real, imag} */,
  {32'hc290754c, 32'hc2d6a36f} /* (16, 13, 25) {real, imag} */,
  {32'hc25d9748, 32'hc123d8e0} /* (16, 13, 24) {real, imag} */,
  {32'h41d8b0b2, 32'h4200f784} /* (16, 13, 23) {real, imag} */,
  {32'h42507656, 32'hbf6cd4b0} /* (16, 13, 22) {real, imag} */,
  {32'h4013f4c4, 32'h42597132} /* (16, 13, 21) {real, imag} */,
  {32'h423e83fc, 32'hc1dbba6e} /* (16, 13, 20) {real, imag} */,
  {32'h41288294, 32'hbff536bc} /* (16, 13, 19) {real, imag} */,
  {32'hc23e86c2, 32'h4290dd4f} /* (16, 13, 18) {real, imag} */,
  {32'hc254d5d6, 32'hc1914caa} /* (16, 13, 17) {real, imag} */,
  {32'hc2097b90, 32'h00000000} /* (16, 13, 16) {real, imag} */,
  {32'hc254d5d6, 32'h41914caa} /* (16, 13, 15) {real, imag} */,
  {32'hc23e86c2, 32'hc290dd4f} /* (16, 13, 14) {real, imag} */,
  {32'h41288294, 32'h3ff536bc} /* (16, 13, 13) {real, imag} */,
  {32'h423e83fc, 32'h41dbba6e} /* (16, 13, 12) {real, imag} */,
  {32'h4013f4c4, 32'hc2597132} /* (16, 13, 11) {real, imag} */,
  {32'h42507656, 32'h3f6cd4b0} /* (16, 13, 10) {real, imag} */,
  {32'h41d8b0b2, 32'hc200f784} /* (16, 13, 9) {real, imag} */,
  {32'hc25d9748, 32'h4123d8e0} /* (16, 13, 8) {real, imag} */,
  {32'hc290754c, 32'h42d6a36f} /* (16, 13, 7) {real, imag} */,
  {32'hc2b31e6e, 32'h41d655fa} /* (16, 13, 6) {real, imag} */,
  {32'hc345b854, 32'hc200665c} /* (16, 13, 5) {real, imag} */,
  {32'h42e219a8, 32'hc2c0a6aa} /* (16, 13, 4) {real, imag} */,
  {32'hc2537f90, 32'hc2418122} /* (16, 13, 3) {real, imag} */,
  {32'hc3a33508, 32'hc2a01623} /* (16, 13, 2) {real, imag} */,
  {32'h442bb184, 32'hc3455032} /* (16, 13, 1) {real, imag} */,
  {32'h444010bd, 32'h00000000} /* (16, 13, 0) {real, imag} */,
  {32'h44182680, 32'h431bb5c3} /* (16, 12, 31) {real, imag} */,
  {32'hc3c138bc, 32'h42c46d1f} /* (16, 12, 30) {real, imag} */,
  {32'h42af6a29, 32'h429b1f3f} /* (16, 12, 29) {real, imag} */,
  {32'h40eaa480, 32'h42c22e89} /* (16, 12, 28) {real, imag} */,
  {32'hc2a919a2, 32'h42a8ce1f} /* (16, 12, 27) {real, imag} */,
  {32'h425ee502, 32'h425a9ee2} /* (16, 12, 26) {real, imag} */,
  {32'hc2acd686, 32'hc18db5b2} /* (16, 12, 25) {real, imag} */,
  {32'hc22eeee0, 32'h430b3c16} /* (16, 12, 24) {real, imag} */,
  {32'h417a0858, 32'hc2b155b2} /* (16, 12, 23) {real, imag} */,
  {32'h415830b0, 32'h423e0582} /* (16, 12, 22) {real, imag} */,
  {32'h404cf240, 32'h42095291} /* (16, 12, 21) {real, imag} */,
  {32'h419c35e4, 32'hc223c2e1} /* (16, 12, 20) {real, imag} */,
  {32'hc2193a68, 32'hc21b45b4} /* (16, 12, 19) {real, imag} */,
  {32'hbe723bc0, 32'hc2a20248} /* (16, 12, 18) {real, imag} */,
  {32'h425102ed, 32'hc2810332} /* (16, 12, 17) {real, imag} */,
  {32'hc22d94bc, 32'h00000000} /* (16, 12, 16) {real, imag} */,
  {32'h425102ed, 32'h42810332} /* (16, 12, 15) {real, imag} */,
  {32'hbe723bc0, 32'h42a20248} /* (16, 12, 14) {real, imag} */,
  {32'hc2193a68, 32'h421b45b4} /* (16, 12, 13) {real, imag} */,
  {32'h419c35e4, 32'h4223c2e1} /* (16, 12, 12) {real, imag} */,
  {32'h404cf240, 32'hc2095291} /* (16, 12, 11) {real, imag} */,
  {32'h415830b0, 32'hc23e0582} /* (16, 12, 10) {real, imag} */,
  {32'h417a0858, 32'h42b155b2} /* (16, 12, 9) {real, imag} */,
  {32'hc22eeee0, 32'hc30b3c16} /* (16, 12, 8) {real, imag} */,
  {32'hc2acd686, 32'h418db5b2} /* (16, 12, 7) {real, imag} */,
  {32'h425ee502, 32'hc25a9ee2} /* (16, 12, 6) {real, imag} */,
  {32'hc2a919a2, 32'hc2a8ce1f} /* (16, 12, 5) {real, imag} */,
  {32'h40eaa480, 32'hc2c22e89} /* (16, 12, 4) {real, imag} */,
  {32'h42af6a29, 32'hc29b1f3f} /* (16, 12, 3) {real, imag} */,
  {32'hc3c138bc, 32'hc2c46d1f} /* (16, 12, 2) {real, imag} */,
  {32'h44182680, 32'hc31bb5c3} /* (16, 12, 1) {real, imag} */,
  {32'h446a6db6, 32'h00000000} /* (16, 12, 0) {real, imag} */,
  {32'h43a17cfa, 32'h43a1fc44} /* (16, 11, 31) {real, imag} */,
  {32'hc37190ea, 32'h43090805} /* (16, 11, 30) {real, imag} */,
  {32'h424eff25, 32'hc28bf662} /* (16, 11, 29) {real, imag} */,
  {32'hc1feeaad, 32'hc30c9656} /* (16, 11, 28) {real, imag} */,
  {32'hc2989473, 32'h4213c534} /* (16, 11, 27) {real, imag} */,
  {32'h42c01bde, 32'h42a4039e} /* (16, 11, 26) {real, imag} */,
  {32'h422f02bf, 32'hc2ddd486} /* (16, 11, 25) {real, imag} */,
  {32'h41e3b18f, 32'h4312878f} /* (16, 11, 24) {real, imag} */,
  {32'hc1e89969, 32'hc25ee5e2} /* (16, 11, 23) {real, imag} */,
  {32'hc31c6f16, 32'h41a9e8ae} /* (16, 11, 22) {real, imag} */,
  {32'h424a1391, 32'h3fef7a08} /* (16, 11, 21) {real, imag} */,
  {32'h42fa79a8, 32'h425018a7} /* (16, 11, 20) {real, imag} */,
  {32'hc210d0fd, 32'h4272a1bd} /* (16, 11, 19) {real, imag} */,
  {32'h3febc318, 32'h41f4993e} /* (16, 11, 18) {real, imag} */,
  {32'h4248e594, 32'hc23604cb} /* (16, 11, 17) {real, imag} */,
  {32'h42a1be04, 32'h00000000} /* (16, 11, 16) {real, imag} */,
  {32'h4248e594, 32'h423604cb} /* (16, 11, 15) {real, imag} */,
  {32'h3febc318, 32'hc1f4993e} /* (16, 11, 14) {real, imag} */,
  {32'hc210d0fd, 32'hc272a1bd} /* (16, 11, 13) {real, imag} */,
  {32'h42fa79a8, 32'hc25018a7} /* (16, 11, 12) {real, imag} */,
  {32'h424a1391, 32'hbfef7a08} /* (16, 11, 11) {real, imag} */,
  {32'hc31c6f16, 32'hc1a9e8ae} /* (16, 11, 10) {real, imag} */,
  {32'hc1e89969, 32'h425ee5e2} /* (16, 11, 9) {real, imag} */,
  {32'h41e3b18f, 32'hc312878f} /* (16, 11, 8) {real, imag} */,
  {32'h422f02bf, 32'h42ddd486} /* (16, 11, 7) {real, imag} */,
  {32'h42c01bde, 32'hc2a4039e} /* (16, 11, 6) {real, imag} */,
  {32'hc2989473, 32'hc213c534} /* (16, 11, 5) {real, imag} */,
  {32'hc1feeaad, 32'h430c9656} /* (16, 11, 4) {real, imag} */,
  {32'h424eff25, 32'h428bf662} /* (16, 11, 3) {real, imag} */,
  {32'hc37190ea, 32'hc3090805} /* (16, 11, 2) {real, imag} */,
  {32'h43a17cfa, 32'hc3a1fc44} /* (16, 11, 1) {real, imag} */,
  {32'h445d321b, 32'h00000000} /* (16, 11, 0) {real, imag} */,
  {32'hc3b2aedd, 32'h43b4bc28} /* (16, 10, 31) {real, imag} */,
  {32'h43622238, 32'h42ba361e} /* (16, 10, 30) {real, imag} */,
  {32'hc29f11c0, 32'hc233fbe2} /* (16, 10, 29) {real, imag} */,
  {32'hc1d461c0, 32'hc280ce1c} /* (16, 10, 28) {real, imag} */,
  {32'hc1a99512, 32'hc2062650} /* (16, 10, 27) {real, imag} */,
  {32'hc207671a, 32'h421f1426} /* (16, 10, 26) {real, imag} */,
  {32'hc10f0cfe, 32'h42daf137} /* (16, 10, 25) {real, imag} */,
  {32'h3fa27ce0, 32'h40e06f80} /* (16, 10, 24) {real, imag} */,
  {32'hbefcb8c0, 32'h428b68fe} /* (16, 10, 23) {real, imag} */,
  {32'h42284e9c, 32'hc2bbe15c} /* (16, 10, 22) {real, imag} */,
  {32'h421f7240, 32'hbf80bb20} /* (16, 10, 21) {real, imag} */,
  {32'h41dbcec6, 32'hc16c1ba8} /* (16, 10, 20) {real, imag} */,
  {32'h428c4b25, 32'h42c589bf} /* (16, 10, 19) {real, imag} */,
  {32'hc1f164fe, 32'hc21d4769} /* (16, 10, 18) {real, imag} */,
  {32'h420139ac, 32'hc20df39a} /* (16, 10, 17) {real, imag} */,
  {32'h423397c3, 32'h00000000} /* (16, 10, 16) {real, imag} */,
  {32'h420139ac, 32'h420df39a} /* (16, 10, 15) {real, imag} */,
  {32'hc1f164fe, 32'h421d4769} /* (16, 10, 14) {real, imag} */,
  {32'h428c4b25, 32'hc2c589bf} /* (16, 10, 13) {real, imag} */,
  {32'h41dbcec6, 32'h416c1ba8} /* (16, 10, 12) {real, imag} */,
  {32'h421f7240, 32'h3f80bb20} /* (16, 10, 11) {real, imag} */,
  {32'h42284e9c, 32'h42bbe15c} /* (16, 10, 10) {real, imag} */,
  {32'hbefcb8c0, 32'hc28b68fe} /* (16, 10, 9) {real, imag} */,
  {32'h3fa27ce0, 32'hc0e06f80} /* (16, 10, 8) {real, imag} */,
  {32'hc10f0cfe, 32'hc2daf137} /* (16, 10, 7) {real, imag} */,
  {32'hc207671a, 32'hc21f1426} /* (16, 10, 6) {real, imag} */,
  {32'hc1a99512, 32'h42062650} /* (16, 10, 5) {real, imag} */,
  {32'hc1d461c0, 32'h4280ce1c} /* (16, 10, 4) {real, imag} */,
  {32'hc29f11c0, 32'h4233fbe2} /* (16, 10, 3) {real, imag} */,
  {32'h43622238, 32'hc2ba361e} /* (16, 10, 2) {real, imag} */,
  {32'hc3b2aedd, 32'hc3b4bc28} /* (16, 10, 1) {real, imag} */,
  {32'h438b907e, 32'h00000000} /* (16, 10, 0) {real, imag} */,
  {32'hc4511574, 32'h439baf47} /* (16, 9, 31) {real, imag} */,
  {32'h43da9751, 32'hc09cfdbc} /* (16, 9, 30) {real, imag} */,
  {32'hc3188913, 32'h42847bed} /* (16, 9, 29) {real, imag} */,
  {32'h40a63480, 32'h42358a78} /* (16, 9, 28) {real, imag} */,
  {32'h4275dded, 32'hc195f2d8} /* (16, 9, 27) {real, imag} */,
  {32'h4185f858, 32'hc1020ea2} /* (16, 9, 26) {real, imag} */,
  {32'hc2f702f6, 32'h42f831da} /* (16, 9, 25) {real, imag} */,
  {32'h42337d25, 32'hc22dbf18} /* (16, 9, 24) {real, imag} */,
  {32'h42a70b15, 32'hc221fce3} /* (16, 9, 23) {real, imag} */,
  {32'h4241ff82, 32'hc189e844} /* (16, 9, 22) {real, imag} */,
  {32'h4299a9b1, 32'h4105c4b8} /* (16, 9, 21) {real, imag} */,
  {32'hc28cdd62, 32'hc19cdbbc} /* (16, 9, 20) {real, imag} */,
  {32'hc2c07719, 32'hc1cc452a} /* (16, 9, 19) {real, imag} */,
  {32'hc28f0ce7, 32'h41a12a7c} /* (16, 9, 18) {real, imag} */,
  {32'h421f2f44, 32'h4195b1ce} /* (16, 9, 17) {real, imag} */,
  {32'hc1b93228, 32'h00000000} /* (16, 9, 16) {real, imag} */,
  {32'h421f2f44, 32'hc195b1ce} /* (16, 9, 15) {real, imag} */,
  {32'hc28f0ce7, 32'hc1a12a7c} /* (16, 9, 14) {real, imag} */,
  {32'hc2c07719, 32'h41cc452a} /* (16, 9, 13) {real, imag} */,
  {32'hc28cdd62, 32'h419cdbbc} /* (16, 9, 12) {real, imag} */,
  {32'h4299a9b1, 32'hc105c4b8} /* (16, 9, 11) {real, imag} */,
  {32'h4241ff82, 32'h4189e844} /* (16, 9, 10) {real, imag} */,
  {32'h42a70b15, 32'h4221fce3} /* (16, 9, 9) {real, imag} */,
  {32'h42337d25, 32'h422dbf18} /* (16, 9, 8) {real, imag} */,
  {32'hc2f702f6, 32'hc2f831da} /* (16, 9, 7) {real, imag} */,
  {32'h4185f858, 32'h41020ea2} /* (16, 9, 6) {real, imag} */,
  {32'h4275dded, 32'h4195f2d8} /* (16, 9, 5) {real, imag} */,
  {32'h40a63480, 32'hc2358a78} /* (16, 9, 4) {real, imag} */,
  {32'hc3188913, 32'hc2847bed} /* (16, 9, 3) {real, imag} */,
  {32'h43da9751, 32'h409cfdbc} /* (16, 9, 2) {real, imag} */,
  {32'hc4511574, 32'hc39baf47} /* (16, 9, 1) {real, imag} */,
  {32'hc309ca3c, 32'h00000000} /* (16, 9, 0) {real, imag} */,
  {32'hc483e942, 32'h43aa6950} /* (16, 8, 31) {real, imag} */,
  {32'h43accb02, 32'hc3095eae} /* (16, 8, 30) {real, imag} */,
  {32'hc380556a, 32'hc1278910} /* (16, 8, 29) {real, imag} */,
  {32'hc28e7eb8, 32'h41643790} /* (16, 8, 28) {real, imag} */,
  {32'hc0f4ad80, 32'hc104d8f0} /* (16, 8, 27) {real, imag} */,
  {32'hc2fec4fe, 32'h4216cfb8} /* (16, 8, 26) {real, imag} */,
  {32'hc2a40c96, 32'hc2aacc40} /* (16, 8, 25) {real, imag} */,
  {32'h4227b3b3, 32'hc2fe5492} /* (16, 8, 24) {real, imag} */,
  {32'hc1c82bd0, 32'hc2bc5081} /* (16, 8, 23) {real, imag} */,
  {32'hc0e3d7d0, 32'hc24c51ec} /* (16, 8, 22) {real, imag} */,
  {32'hc2d88d8b, 32'hc1d8a415} /* (16, 8, 21) {real, imag} */,
  {32'h426e0350, 32'h4292ef16} /* (16, 8, 20) {real, imag} */,
  {32'hc2b21308, 32'hc246daca} /* (16, 8, 19) {real, imag} */,
  {32'hc2173112, 32'h420030bd} /* (16, 8, 18) {real, imag} */,
  {32'hc0413784, 32'hc22969a7} /* (16, 8, 17) {real, imag} */,
  {32'h42048f90, 32'h00000000} /* (16, 8, 16) {real, imag} */,
  {32'hc0413784, 32'h422969a7} /* (16, 8, 15) {real, imag} */,
  {32'hc2173112, 32'hc20030bd} /* (16, 8, 14) {real, imag} */,
  {32'hc2b21308, 32'h4246daca} /* (16, 8, 13) {real, imag} */,
  {32'h426e0350, 32'hc292ef16} /* (16, 8, 12) {real, imag} */,
  {32'hc2d88d8b, 32'h41d8a415} /* (16, 8, 11) {real, imag} */,
  {32'hc0e3d7d0, 32'h424c51ec} /* (16, 8, 10) {real, imag} */,
  {32'hc1c82bd0, 32'h42bc5081} /* (16, 8, 9) {real, imag} */,
  {32'h4227b3b3, 32'h42fe5492} /* (16, 8, 8) {real, imag} */,
  {32'hc2a40c96, 32'h42aacc40} /* (16, 8, 7) {real, imag} */,
  {32'hc2fec4fe, 32'hc216cfb8} /* (16, 8, 6) {real, imag} */,
  {32'hc0f4ad80, 32'h4104d8f0} /* (16, 8, 5) {real, imag} */,
  {32'hc28e7eb8, 32'hc1643790} /* (16, 8, 4) {real, imag} */,
  {32'hc380556a, 32'h41278910} /* (16, 8, 3) {real, imag} */,
  {32'h43accb02, 32'h43095eae} /* (16, 8, 2) {real, imag} */,
  {32'hc483e942, 32'hc3aa6950} /* (16, 8, 1) {real, imag} */,
  {32'hc3a6b5d9, 32'h00000000} /* (16, 8, 0) {real, imag} */,
  {32'hc486f407, 32'h43f0f183} /* (16, 7, 31) {real, imag} */,
  {32'h438b976d, 32'hc3690d8a} /* (16, 7, 30) {real, imag} */,
  {32'hc2a04ad0, 32'h4218221a} /* (16, 7, 29) {real, imag} */,
  {32'hc2c399c1, 32'hc1b4fd38} /* (16, 7, 28) {real, imag} */,
  {32'h42bff836, 32'hc219e48c} /* (16, 7, 27) {real, imag} */,
  {32'hc20c1c7c, 32'h431f75bf} /* (16, 7, 26) {real, imag} */,
  {32'hc1114edc, 32'hc1ec2e3d} /* (16, 7, 25) {real, imag} */,
  {32'h413cd7a0, 32'hc22947b4} /* (16, 7, 24) {real, imag} */,
  {32'h42494c98, 32'hc273e237} /* (16, 7, 23) {real, imag} */,
  {32'hc186d190, 32'h43025994} /* (16, 7, 22) {real, imag} */,
  {32'h42174173, 32'hc3206349} /* (16, 7, 21) {real, imag} */,
  {32'h42ed9cf8, 32'h41bcfd29} /* (16, 7, 20) {real, imag} */,
  {32'hc19a41b9, 32'hc17fdc7e} /* (16, 7, 19) {real, imag} */,
  {32'h41de0806, 32'h4196ab49} /* (16, 7, 18) {real, imag} */,
  {32'h4192a61e, 32'h42a5bd02} /* (16, 7, 17) {real, imag} */,
  {32'hc310dd18, 32'h00000000} /* (16, 7, 16) {real, imag} */,
  {32'h4192a61e, 32'hc2a5bd02} /* (16, 7, 15) {real, imag} */,
  {32'h41de0806, 32'hc196ab49} /* (16, 7, 14) {real, imag} */,
  {32'hc19a41b9, 32'h417fdc7e} /* (16, 7, 13) {real, imag} */,
  {32'h42ed9cf8, 32'hc1bcfd29} /* (16, 7, 12) {real, imag} */,
  {32'h42174173, 32'h43206349} /* (16, 7, 11) {real, imag} */,
  {32'hc186d190, 32'hc3025994} /* (16, 7, 10) {real, imag} */,
  {32'h42494c98, 32'h4273e237} /* (16, 7, 9) {real, imag} */,
  {32'h413cd7a0, 32'h422947b4} /* (16, 7, 8) {real, imag} */,
  {32'hc1114edc, 32'h41ec2e3d} /* (16, 7, 7) {real, imag} */,
  {32'hc20c1c7c, 32'hc31f75bf} /* (16, 7, 6) {real, imag} */,
  {32'h42bff836, 32'h4219e48c} /* (16, 7, 5) {real, imag} */,
  {32'hc2c399c1, 32'h41b4fd38} /* (16, 7, 4) {real, imag} */,
  {32'hc2a04ad0, 32'hc218221a} /* (16, 7, 3) {real, imag} */,
  {32'h438b976d, 32'h43690d8a} /* (16, 7, 2) {real, imag} */,
  {32'hc486f407, 32'hc3f0f183} /* (16, 7, 1) {real, imag} */,
  {32'hc431f69c, 32'h00000000} /* (16, 7, 0) {real, imag} */,
  {32'hc48a543d, 32'h44080290} /* (16, 6, 31) {real, imag} */,
  {32'h4360c70e, 32'hc331368c} /* (16, 6, 30) {real, imag} */,
  {32'hc2c6d490, 32'hc1113d08} /* (16, 6, 29) {real, imag} */,
  {32'hc251cabc, 32'hc20fc19d} /* (16, 6, 28) {real, imag} */,
  {32'h42a95600, 32'hc2ee5d04} /* (16, 6, 27) {real, imag} */,
  {32'h420ce9c0, 32'hc1bf2ace} /* (16, 6, 26) {real, imag} */,
  {32'h41c2013d, 32'h402ee7b8} /* (16, 6, 25) {real, imag} */,
  {32'h423a49ae, 32'hc31090c5} /* (16, 6, 24) {real, imag} */,
  {32'hc03bbb20, 32'hc1911724} /* (16, 6, 23) {real, imag} */,
  {32'hc220a72f, 32'h42b898d1} /* (16, 6, 22) {real, imag} */,
  {32'hc28f495a, 32'hc223afe5} /* (16, 6, 21) {real, imag} */,
  {32'h42d50212, 32'hc22373aa} /* (16, 6, 20) {real, imag} */,
  {32'h42761dc9, 32'h4265719a} /* (16, 6, 19) {real, imag} */,
  {32'h414f61d5, 32'hc24bdab8} /* (16, 6, 18) {real, imag} */,
  {32'h4234a941, 32'h41ba5d78} /* (16, 6, 17) {real, imag} */,
  {32'hc0e0c320, 32'h00000000} /* (16, 6, 16) {real, imag} */,
  {32'h4234a941, 32'hc1ba5d78} /* (16, 6, 15) {real, imag} */,
  {32'h414f61d5, 32'h424bdab8} /* (16, 6, 14) {real, imag} */,
  {32'h42761dc9, 32'hc265719a} /* (16, 6, 13) {real, imag} */,
  {32'h42d50212, 32'h422373aa} /* (16, 6, 12) {real, imag} */,
  {32'hc28f495a, 32'h4223afe5} /* (16, 6, 11) {real, imag} */,
  {32'hc220a72f, 32'hc2b898d1} /* (16, 6, 10) {real, imag} */,
  {32'hc03bbb20, 32'h41911724} /* (16, 6, 9) {real, imag} */,
  {32'h423a49ae, 32'h431090c5} /* (16, 6, 8) {real, imag} */,
  {32'h41c2013d, 32'hc02ee7b8} /* (16, 6, 7) {real, imag} */,
  {32'h420ce9c0, 32'h41bf2ace} /* (16, 6, 6) {real, imag} */,
  {32'h42a95600, 32'h42ee5d04} /* (16, 6, 5) {real, imag} */,
  {32'hc251cabc, 32'h420fc19d} /* (16, 6, 4) {real, imag} */,
  {32'hc2c6d490, 32'h41113d08} /* (16, 6, 3) {real, imag} */,
  {32'h4360c70e, 32'h4331368c} /* (16, 6, 2) {real, imag} */,
  {32'hc48a543d, 32'hc4080290} /* (16, 6, 1) {real, imag} */,
  {32'hc43a5c44, 32'h00000000} /* (16, 6, 0) {real, imag} */,
  {32'hc47f8c66, 32'h44456861} /* (16, 5, 31) {real, imag} */,
  {32'hc2b7241e, 32'hc38849ac} /* (16, 5, 30) {real, imag} */,
  {32'hc2b138b0, 32'hc2940ea4} /* (16, 5, 29) {real, imag} */,
  {32'h42f29c62, 32'hc2c99de0} /* (16, 5, 28) {real, imag} */,
  {32'h432c694c, 32'hc19d63ce} /* (16, 5, 27) {real, imag} */,
  {32'hc200d67e, 32'hc299e81b} /* (16, 5, 26) {real, imag} */,
  {32'h43076c07, 32'h420ec2b2} /* (16, 5, 25) {real, imag} */,
  {32'h429afc66, 32'hc23254f6} /* (16, 5, 24) {real, imag} */,
  {32'h41b4f82b, 32'hc19b306d} /* (16, 5, 23) {real, imag} */,
  {32'h425484e4, 32'hc248d8dc} /* (16, 5, 22) {real, imag} */,
  {32'hc29088aa, 32'hbf7dd180} /* (16, 5, 21) {real, imag} */,
  {32'hbfba1ab8, 32'h42714521} /* (16, 5, 20) {real, imag} */,
  {32'h425be344, 32'hc27c2070} /* (16, 5, 19) {real, imag} */,
  {32'hc2010bef, 32'hc1d85924} /* (16, 5, 18) {real, imag} */,
  {32'hc26e16ac, 32'hc26d7ec4} /* (16, 5, 17) {real, imag} */,
  {32'hc1178f7b, 32'h00000000} /* (16, 5, 16) {real, imag} */,
  {32'hc26e16ac, 32'h426d7ec4} /* (16, 5, 15) {real, imag} */,
  {32'hc2010bef, 32'h41d85924} /* (16, 5, 14) {real, imag} */,
  {32'h425be344, 32'h427c2070} /* (16, 5, 13) {real, imag} */,
  {32'hbfba1ab8, 32'hc2714521} /* (16, 5, 12) {real, imag} */,
  {32'hc29088aa, 32'h3f7dd180} /* (16, 5, 11) {real, imag} */,
  {32'h425484e4, 32'h4248d8dc} /* (16, 5, 10) {real, imag} */,
  {32'h41b4f82b, 32'h419b306d} /* (16, 5, 9) {real, imag} */,
  {32'h429afc66, 32'h423254f6} /* (16, 5, 8) {real, imag} */,
  {32'h43076c07, 32'hc20ec2b2} /* (16, 5, 7) {real, imag} */,
  {32'hc200d67e, 32'h4299e81b} /* (16, 5, 6) {real, imag} */,
  {32'h432c694c, 32'h419d63ce} /* (16, 5, 5) {real, imag} */,
  {32'h42f29c62, 32'h42c99de0} /* (16, 5, 4) {real, imag} */,
  {32'hc2b138b0, 32'h42940ea4} /* (16, 5, 3) {real, imag} */,
  {32'hc2b7241e, 32'h438849ac} /* (16, 5, 2) {real, imag} */,
  {32'hc47f8c66, 32'hc4456861} /* (16, 5, 1) {real, imag} */,
  {32'hc4462805, 32'h00000000} /* (16, 5, 0) {real, imag} */,
  {32'hc4333586, 32'h4469f7ac} /* (16, 4, 31) {real, imag} */,
  {32'hc3c84819, 32'hc3bc9c3d} /* (16, 4, 30) {real, imag} */,
  {32'h41640d8a, 32'h4230bded} /* (16, 4, 29) {real, imag} */,
  {32'h430bfe47, 32'hc33474fa} /* (16, 4, 28) {real, imag} */,
  {32'h4333d1c0, 32'hc1c6ca6d} /* (16, 4, 27) {real, imag} */,
  {32'h4202dbc9, 32'h42bc70d6} /* (16, 4, 26) {real, imag} */,
  {32'h433559ec, 32'hc27cb058} /* (16, 4, 25) {real, imag} */,
  {32'hc319dcc6, 32'h412b15b8} /* (16, 4, 24) {real, imag} */,
  {32'h41059bb8, 32'h41f400c6} /* (16, 4, 23) {real, imag} */,
  {32'hc2fb8e5a, 32'hc2b22f08} /* (16, 4, 22) {real, imag} */,
  {32'h41136ef4, 32'hc24ef644} /* (16, 4, 21) {real, imag} */,
  {32'h42094a65, 32'h42acc0d6} /* (16, 4, 20) {real, imag} */,
  {32'hc2a9ba5b, 32'h41ba4324} /* (16, 4, 19) {real, imag} */,
  {32'hc1ca78e4, 32'h422b9db4} /* (16, 4, 18) {real, imag} */,
  {32'h4037295d, 32'hc0fbf62c} /* (16, 4, 17) {real, imag} */,
  {32'hc2929778, 32'h00000000} /* (16, 4, 16) {real, imag} */,
  {32'h4037295d, 32'h40fbf62c} /* (16, 4, 15) {real, imag} */,
  {32'hc1ca78e4, 32'hc22b9db4} /* (16, 4, 14) {real, imag} */,
  {32'hc2a9ba5b, 32'hc1ba4324} /* (16, 4, 13) {real, imag} */,
  {32'h42094a65, 32'hc2acc0d6} /* (16, 4, 12) {real, imag} */,
  {32'h41136ef4, 32'h424ef644} /* (16, 4, 11) {real, imag} */,
  {32'hc2fb8e5a, 32'h42b22f08} /* (16, 4, 10) {real, imag} */,
  {32'h41059bb8, 32'hc1f400c6} /* (16, 4, 9) {real, imag} */,
  {32'hc319dcc6, 32'hc12b15b8} /* (16, 4, 8) {real, imag} */,
  {32'h433559ec, 32'h427cb058} /* (16, 4, 7) {real, imag} */,
  {32'h4202dbc9, 32'hc2bc70d6} /* (16, 4, 6) {real, imag} */,
  {32'h4333d1c0, 32'h41c6ca6d} /* (16, 4, 5) {real, imag} */,
  {32'h430bfe47, 32'h433474fa} /* (16, 4, 4) {real, imag} */,
  {32'h41640d8a, 32'hc230bded} /* (16, 4, 3) {real, imag} */,
  {32'hc3c84819, 32'h43bc9c3d} /* (16, 4, 2) {real, imag} */,
  {32'hc4333586, 32'hc469f7ac} /* (16, 4, 1) {real, imag} */,
  {32'hc43c66b5, 32'h00000000} /* (16, 4, 0) {real, imag} */,
  {32'hc41443ea, 32'h4477b4e0} /* (16, 3, 31) {real, imag} */,
  {32'hc375c364, 32'hc3abea61} /* (16, 3, 30) {real, imag} */,
  {32'h422b77ec, 32'h42f9ea53} /* (16, 3, 29) {real, imag} */,
  {32'h42502202, 32'hc26f1d7c} /* (16, 3, 28) {real, imag} */,
  {32'h42cc67bc, 32'h43044137} /* (16, 3, 27) {real, imag} */,
  {32'h41aa4c0c, 32'hc18a7228} /* (16, 3, 26) {real, imag} */,
  {32'h4233f1d4, 32'h428d2366} /* (16, 3, 25) {real, imag} */,
  {32'h3f946210, 32'hc2c47998} /* (16, 3, 24) {real, imag} */,
  {32'h41c0a94a, 32'hc21857da} /* (16, 3, 23) {real, imag} */,
  {32'h41aa3508, 32'hc23b6d42} /* (16, 3, 22) {real, imag} */,
  {32'h41a07df0, 32'hc2baebb5} /* (16, 3, 21) {real, imag} */,
  {32'h401a99e0, 32'h42af9026} /* (16, 3, 20) {real, imag} */,
  {32'hc27aa943, 32'h417bcf4a} /* (16, 3, 19) {real, imag} */,
  {32'hc22304ce, 32'h4267bfca} /* (16, 3, 18) {real, imag} */,
  {32'h4217228e, 32'hc27aeb6c} /* (16, 3, 17) {real, imag} */,
  {32'hc0d5e44e, 32'h00000000} /* (16, 3, 16) {real, imag} */,
  {32'h4217228e, 32'h427aeb6c} /* (16, 3, 15) {real, imag} */,
  {32'hc22304ce, 32'hc267bfca} /* (16, 3, 14) {real, imag} */,
  {32'hc27aa943, 32'hc17bcf4a} /* (16, 3, 13) {real, imag} */,
  {32'h401a99e0, 32'hc2af9026} /* (16, 3, 12) {real, imag} */,
  {32'h41a07df0, 32'h42baebb5} /* (16, 3, 11) {real, imag} */,
  {32'h41aa3508, 32'h423b6d42} /* (16, 3, 10) {real, imag} */,
  {32'h41c0a94a, 32'h421857da} /* (16, 3, 9) {real, imag} */,
  {32'h3f946210, 32'h42c47998} /* (16, 3, 8) {real, imag} */,
  {32'h4233f1d4, 32'hc28d2366} /* (16, 3, 7) {real, imag} */,
  {32'h41aa4c0c, 32'h418a7228} /* (16, 3, 6) {real, imag} */,
  {32'h42cc67bc, 32'hc3044137} /* (16, 3, 5) {real, imag} */,
  {32'h42502202, 32'h426f1d7c} /* (16, 3, 4) {real, imag} */,
  {32'h422b77ec, 32'hc2f9ea53} /* (16, 3, 3) {real, imag} */,
  {32'hc375c364, 32'h43abea61} /* (16, 3, 2) {real, imag} */,
  {32'hc41443ea, 32'hc477b4e0} /* (16, 3, 1) {real, imag} */,
  {32'hc43aa1b4, 32'h00000000} /* (16, 3, 0) {real, imag} */,
  {32'hc4212180, 32'h44731b40} /* (16, 2, 31) {real, imag} */,
  {32'hc31e6b83, 32'hc3eabbf9} /* (16, 2, 30) {real, imag} */,
  {32'h431622a4, 32'h4297cd92} /* (16, 2, 29) {real, imag} */,
  {32'h41c9a9ed, 32'hc36909f4} /* (16, 2, 28) {real, imag} */,
  {32'hc14cd510, 32'h42eb3a54} /* (16, 2, 27) {real, imag} */,
  {32'hc1aaf558, 32'hc28ed7ea} /* (16, 2, 26) {real, imag} */,
  {32'h422749ab, 32'h4213a2e4} /* (16, 2, 25) {real, imag} */,
  {32'h42dcd4a4, 32'hc22ae740} /* (16, 2, 24) {real, imag} */,
  {32'hc2b6cda1, 32'h41594ca3} /* (16, 2, 23) {real, imag} */,
  {32'h42a2a951, 32'h41e6f7ad} /* (16, 2, 22) {real, imag} */,
  {32'hc1eef948, 32'h421eb472} /* (16, 2, 21) {real, imag} */,
  {32'h411ecd3a, 32'h416a833a} /* (16, 2, 20) {real, imag} */,
  {32'h41e715fc, 32'h3ff35fd0} /* (16, 2, 19) {real, imag} */,
  {32'h419649b0, 32'hc206fb3a} /* (16, 2, 18) {real, imag} */,
  {32'hc264abe9, 32'h42085c12} /* (16, 2, 17) {real, imag} */,
  {32'hc0d2f05c, 32'h00000000} /* (16, 2, 16) {real, imag} */,
  {32'hc264abe9, 32'hc2085c12} /* (16, 2, 15) {real, imag} */,
  {32'h419649b0, 32'h4206fb3a} /* (16, 2, 14) {real, imag} */,
  {32'h41e715fc, 32'hbff35fd0} /* (16, 2, 13) {real, imag} */,
  {32'h411ecd3a, 32'hc16a833a} /* (16, 2, 12) {real, imag} */,
  {32'hc1eef948, 32'hc21eb472} /* (16, 2, 11) {real, imag} */,
  {32'h42a2a951, 32'hc1e6f7ad} /* (16, 2, 10) {real, imag} */,
  {32'hc2b6cda1, 32'hc1594ca3} /* (16, 2, 9) {real, imag} */,
  {32'h42dcd4a4, 32'h422ae740} /* (16, 2, 8) {real, imag} */,
  {32'h422749ab, 32'hc213a2e4} /* (16, 2, 7) {real, imag} */,
  {32'hc1aaf558, 32'h428ed7ea} /* (16, 2, 6) {real, imag} */,
  {32'hc14cd510, 32'hc2eb3a54} /* (16, 2, 5) {real, imag} */,
  {32'h41c9a9ed, 32'h436909f4} /* (16, 2, 4) {real, imag} */,
  {32'h431622a4, 32'hc297cd92} /* (16, 2, 3) {real, imag} */,
  {32'hc31e6b83, 32'h43eabbf9} /* (16, 2, 2) {real, imag} */,
  {32'hc4212180, 32'hc4731b40} /* (16, 2, 1) {real, imag} */,
  {32'hc451706c, 32'h00000000} /* (16, 2, 0) {real, imag} */,
  {32'hc4323fe7, 32'h44489173} /* (16, 1, 31) {real, imag} */,
  {32'hc2481eb0, 32'hc3e22563} /* (16, 1, 30) {real, imag} */,
  {32'h42ca7525, 32'h43046cf0} /* (16, 1, 29) {real, imag} */,
  {32'h41076248, 32'hc3045d46} /* (16, 1, 28) {real, imag} */,
  {32'h428f581b, 32'h423bb758} /* (16, 1, 27) {real, imag} */,
  {32'h40d2e0f8, 32'hc26d0b3b} /* (16, 1, 26) {real, imag} */,
  {32'hc226c86d, 32'hc20df0f5} /* (16, 1, 25) {real, imag} */,
  {32'h40b6a8d4, 32'hc1950d0b} /* (16, 1, 24) {real, imag} */,
  {32'hc30a9e65, 32'h4222cb54} /* (16, 1, 23) {real, imag} */,
  {32'hc1c448a2, 32'h41a6780b} /* (16, 1, 22) {real, imag} */,
  {32'h426264ce, 32'hc225511c} /* (16, 1, 21) {real, imag} */,
  {32'hc17209a3, 32'hc2902c57} /* (16, 1, 20) {real, imag} */,
  {32'h4202d6e0, 32'h419fcc30} /* (16, 1, 19) {real, imag} */,
  {32'hc1edd279, 32'hc09abe28} /* (16, 1, 18) {real, imag} */,
  {32'hc2b94654, 32'hc2ec1208} /* (16, 1, 17) {real, imag} */,
  {32'hc288ed0c, 32'h00000000} /* (16, 1, 16) {real, imag} */,
  {32'hc2b94654, 32'h42ec1208} /* (16, 1, 15) {real, imag} */,
  {32'hc1edd279, 32'h409abe28} /* (16, 1, 14) {real, imag} */,
  {32'h4202d6e0, 32'hc19fcc30} /* (16, 1, 13) {real, imag} */,
  {32'hc17209a3, 32'h42902c57} /* (16, 1, 12) {real, imag} */,
  {32'h426264ce, 32'h4225511c} /* (16, 1, 11) {real, imag} */,
  {32'hc1c448a2, 32'hc1a6780b} /* (16, 1, 10) {real, imag} */,
  {32'hc30a9e65, 32'hc222cb54} /* (16, 1, 9) {real, imag} */,
  {32'h40b6a8d4, 32'h41950d0b} /* (16, 1, 8) {real, imag} */,
  {32'hc226c86d, 32'h420df0f5} /* (16, 1, 7) {real, imag} */,
  {32'h40d2e0f8, 32'h426d0b3b} /* (16, 1, 6) {real, imag} */,
  {32'h428f581b, 32'hc23bb758} /* (16, 1, 5) {real, imag} */,
  {32'h41076248, 32'h43045d46} /* (16, 1, 4) {real, imag} */,
  {32'h42ca7525, 32'hc3046cf0} /* (16, 1, 3) {real, imag} */,
  {32'hc2481eb0, 32'h43e22563} /* (16, 1, 2) {real, imag} */,
  {32'hc4323fe7, 32'hc4489173} /* (16, 1, 1) {real, imag} */,
  {32'hc468cd18, 32'h00000000} /* (16, 1, 0) {real, imag} */,
  {32'hc42f29f7, 32'h441c302c} /* (16, 0, 31) {real, imag} */,
  {32'h429ab908, 32'hc3b0f986} /* (16, 0, 30) {real, imag} */,
  {32'h423c11c4, 32'h426f9ef0} /* (16, 0, 29) {real, imag} */,
  {32'hc229325a, 32'hc11d8c88} /* (16, 0, 28) {real, imag} */,
  {32'h4231a3cc, 32'h4177aa78} /* (16, 0, 27) {real, imag} */,
  {32'h421bbb52, 32'h4149270c} /* (16, 0, 26) {real, imag} */,
  {32'hc237701e, 32'h4262ada1} /* (16, 0, 25) {real, imag} */,
  {32'hc2240ed6, 32'hc29c7a95} /* (16, 0, 24) {real, imag} */,
  {32'h402118e0, 32'hc20c3e9f} /* (16, 0, 23) {real, imag} */,
  {32'hc1b9ba11, 32'h41947290} /* (16, 0, 22) {real, imag} */,
  {32'h41dce3c4, 32'hc26fb152} /* (16, 0, 21) {real, imag} */,
  {32'hc21a2289, 32'h41f1c670} /* (16, 0, 20) {real, imag} */,
  {32'hc2038c2e, 32'h416fb30a} /* (16, 0, 19) {real, imag} */,
  {32'h411e4ff4, 32'h40b853e4} /* (16, 0, 18) {real, imag} */,
  {32'h412107ee, 32'hc1b18401} /* (16, 0, 17) {real, imag} */,
  {32'hc2bbd458, 32'h00000000} /* (16, 0, 16) {real, imag} */,
  {32'h412107ee, 32'h41b18401} /* (16, 0, 15) {real, imag} */,
  {32'h411e4ff4, 32'hc0b853e4} /* (16, 0, 14) {real, imag} */,
  {32'hc2038c2e, 32'hc16fb30a} /* (16, 0, 13) {real, imag} */,
  {32'hc21a2289, 32'hc1f1c670} /* (16, 0, 12) {real, imag} */,
  {32'h41dce3c4, 32'h426fb152} /* (16, 0, 11) {real, imag} */,
  {32'hc1b9ba11, 32'hc1947290} /* (16, 0, 10) {real, imag} */,
  {32'h402118e0, 32'h420c3e9f} /* (16, 0, 9) {real, imag} */,
  {32'hc2240ed6, 32'h429c7a95} /* (16, 0, 8) {real, imag} */,
  {32'hc237701e, 32'hc262ada1} /* (16, 0, 7) {real, imag} */,
  {32'h421bbb52, 32'hc149270c} /* (16, 0, 6) {real, imag} */,
  {32'h4231a3cc, 32'hc177aa78} /* (16, 0, 5) {real, imag} */,
  {32'hc229325a, 32'h411d8c88} /* (16, 0, 4) {real, imag} */,
  {32'h423c11c4, 32'hc26f9ef0} /* (16, 0, 3) {real, imag} */,
  {32'h429ab908, 32'h43b0f986} /* (16, 0, 2) {real, imag} */,
  {32'hc42f29f7, 32'hc41c302c} /* (16, 0, 1) {real, imag} */,
  {32'hc471de8c, 32'h00000000} /* (16, 0, 0) {real, imag} */,
  {32'h4452e9ad, 32'hc402e741} /* (15, 31, 31) {real, imag} */,
  {32'hc35cdbb9, 32'h43222470} /* (15, 31, 30) {real, imag} */,
  {32'hc1ae8646, 32'h410293b4} /* (15, 31, 29) {real, imag} */,
  {32'h4124effc, 32'hc24286f6} /* (15, 31, 28) {real, imag} */,
  {32'hc2885437, 32'h40b9595c} /* (15, 31, 27) {real, imag} */,
  {32'hc16256fc, 32'h425488e3} /* (15, 31, 26) {real, imag} */,
  {32'h41e4f83d, 32'h4247d328} /* (15, 31, 25) {real, imag} */,
  {32'hc2ef4b80, 32'h41150808} /* (15, 31, 24) {real, imag} */,
  {32'hc2605cae, 32'h4213469e} /* (15, 31, 23) {real, imag} */,
  {32'h41b38bce, 32'hc21e2b9e} /* (15, 31, 22) {real, imag} */,
  {32'h411394b0, 32'h41f50feb} /* (15, 31, 21) {real, imag} */,
  {32'h4247db7d, 32'h41e916d9} /* (15, 31, 20) {real, imag} */,
  {32'hc24d1283, 32'h4236af9e} /* (15, 31, 19) {real, imag} */,
  {32'h41dc577e, 32'hc1cf9428} /* (15, 31, 18) {real, imag} */,
  {32'hc22ec514, 32'hc203e11e} /* (15, 31, 17) {real, imag} */,
  {32'h42017e18, 32'h00000000} /* (15, 31, 16) {real, imag} */,
  {32'hc22ec514, 32'h4203e11e} /* (15, 31, 15) {real, imag} */,
  {32'h41dc577e, 32'h41cf9428} /* (15, 31, 14) {real, imag} */,
  {32'hc24d1283, 32'hc236af9e} /* (15, 31, 13) {real, imag} */,
  {32'h4247db7d, 32'hc1e916d9} /* (15, 31, 12) {real, imag} */,
  {32'h411394b0, 32'hc1f50feb} /* (15, 31, 11) {real, imag} */,
  {32'h41b38bce, 32'h421e2b9e} /* (15, 31, 10) {real, imag} */,
  {32'hc2605cae, 32'hc213469e} /* (15, 31, 9) {real, imag} */,
  {32'hc2ef4b80, 32'hc1150808} /* (15, 31, 8) {real, imag} */,
  {32'h41e4f83d, 32'hc247d328} /* (15, 31, 7) {real, imag} */,
  {32'hc16256fc, 32'hc25488e3} /* (15, 31, 6) {real, imag} */,
  {32'hc2885437, 32'hc0b9595c} /* (15, 31, 5) {real, imag} */,
  {32'h4124effc, 32'h424286f6} /* (15, 31, 4) {real, imag} */,
  {32'hc1ae8646, 32'hc10293b4} /* (15, 31, 3) {real, imag} */,
  {32'hc35cdbb9, 32'hc3222470} /* (15, 31, 2) {real, imag} */,
  {32'h4452e9ad, 32'h4402e741} /* (15, 31, 1) {real, imag} */,
  {32'h4447a1e3, 32'h00000000} /* (15, 31, 0) {real, imag} */,
  {32'h4452e489, 32'hc3d68802} /* (15, 30, 31) {real, imag} */,
  {32'hc3afaaea, 32'h43320c0d} /* (15, 30, 30) {real, imag} */,
  {32'h429356d5, 32'h42ac446a} /* (15, 30, 29) {real, imag} */,
  {32'h42ebead8, 32'hc2c3fb12} /* (15, 30, 28) {real, imag} */,
  {32'h4169c438, 32'h427aa1c8} /* (15, 30, 27) {real, imag} */,
  {32'h42b5bed3, 32'hc0f529e4} /* (15, 30, 26) {real, imag} */,
  {32'h431ea5da, 32'h432e5d56} /* (15, 30, 25) {real, imag} */,
  {32'hc2bc30fc, 32'h422683a0} /* (15, 30, 24) {real, imag} */,
  {32'hc08f8870, 32'h42bc4e8e} /* (15, 30, 23) {real, imag} */,
  {32'hc2941d70, 32'hc1f1b2f4} /* (15, 30, 22) {real, imag} */,
  {32'hc2346182, 32'hc263d68e} /* (15, 30, 21) {real, imag} */,
  {32'h42ad7a51, 32'h42962f4b} /* (15, 30, 20) {real, imag} */,
  {32'h42037776, 32'h4311b916} /* (15, 30, 19) {real, imag} */,
  {32'hc12cd632, 32'h413c53d8} /* (15, 30, 18) {real, imag} */,
  {32'h40c83b76, 32'h4197f926} /* (15, 30, 17) {real, imag} */,
  {32'hc26a68dc, 32'h00000000} /* (15, 30, 16) {real, imag} */,
  {32'h40c83b76, 32'hc197f926} /* (15, 30, 15) {real, imag} */,
  {32'hc12cd632, 32'hc13c53d8} /* (15, 30, 14) {real, imag} */,
  {32'h42037776, 32'hc311b916} /* (15, 30, 13) {real, imag} */,
  {32'h42ad7a51, 32'hc2962f4b} /* (15, 30, 12) {real, imag} */,
  {32'hc2346182, 32'h4263d68e} /* (15, 30, 11) {real, imag} */,
  {32'hc2941d70, 32'h41f1b2f4} /* (15, 30, 10) {real, imag} */,
  {32'hc08f8870, 32'hc2bc4e8e} /* (15, 30, 9) {real, imag} */,
  {32'hc2bc30fc, 32'hc22683a0} /* (15, 30, 8) {real, imag} */,
  {32'h431ea5da, 32'hc32e5d56} /* (15, 30, 7) {real, imag} */,
  {32'h42b5bed3, 32'h40f529e4} /* (15, 30, 6) {real, imag} */,
  {32'h4169c438, 32'hc27aa1c8} /* (15, 30, 5) {real, imag} */,
  {32'h42ebead8, 32'h42c3fb12} /* (15, 30, 4) {real, imag} */,
  {32'h429356d5, 32'hc2ac446a} /* (15, 30, 3) {real, imag} */,
  {32'hc3afaaea, 32'hc3320c0d} /* (15, 30, 2) {real, imag} */,
  {32'h4452e489, 32'h43d68802} /* (15, 30, 1) {real, imag} */,
  {32'h446f2e4e, 32'h00000000} /* (15, 30, 0) {real, imag} */,
  {32'h44219be3, 32'hc3c580ec} /* (15, 29, 31) {real, imag} */,
  {32'hc3e7a030, 32'h42b40424} /* (15, 29, 30) {real, imag} */,
  {32'h4281fea0, 32'h41b511fe} /* (15, 29, 29) {real, imag} */,
  {32'hc28b0580, 32'hc2af756a} /* (15, 29, 28) {real, imag} */,
  {32'h4231fac5, 32'hc0993e60} /* (15, 29, 27) {real, imag} */,
  {32'h430a0b8d, 32'h41ac0c91} /* (15, 29, 26) {real, imag} */,
  {32'h43118b01, 32'hc185ad22} /* (15, 29, 25) {real, imag} */,
  {32'h42514f38, 32'h428c4416} /* (15, 29, 24) {real, imag} */,
  {32'h407e79c0, 32'hc20a505f} /* (15, 29, 23) {real, imag} */,
  {32'hc2c8a1e1, 32'hc1e85d80} /* (15, 29, 22) {real, imag} */,
  {32'hc28b4c81, 32'h4285e3a8} /* (15, 29, 21) {real, imag} */,
  {32'hc1bdf1d8, 32'h417d1fe4} /* (15, 29, 20) {real, imag} */,
  {32'h42b431ca, 32'hc0d4ade8} /* (15, 29, 19) {real, imag} */,
  {32'h4218a650, 32'h421d6c95} /* (15, 29, 18) {real, imag} */,
  {32'h427f7364, 32'h4258fe91} /* (15, 29, 17) {real, imag} */,
  {32'hc2131adf, 32'h00000000} /* (15, 29, 16) {real, imag} */,
  {32'h427f7364, 32'hc258fe91} /* (15, 29, 15) {real, imag} */,
  {32'h4218a650, 32'hc21d6c95} /* (15, 29, 14) {real, imag} */,
  {32'h42b431ca, 32'h40d4ade8} /* (15, 29, 13) {real, imag} */,
  {32'hc1bdf1d8, 32'hc17d1fe4} /* (15, 29, 12) {real, imag} */,
  {32'hc28b4c81, 32'hc285e3a8} /* (15, 29, 11) {real, imag} */,
  {32'hc2c8a1e1, 32'h41e85d80} /* (15, 29, 10) {real, imag} */,
  {32'h407e79c0, 32'h420a505f} /* (15, 29, 9) {real, imag} */,
  {32'h42514f38, 32'hc28c4416} /* (15, 29, 8) {real, imag} */,
  {32'h43118b01, 32'h4185ad22} /* (15, 29, 7) {real, imag} */,
  {32'h430a0b8d, 32'hc1ac0c91} /* (15, 29, 6) {real, imag} */,
  {32'h4231fac5, 32'h40993e60} /* (15, 29, 5) {real, imag} */,
  {32'hc28b0580, 32'h42af756a} /* (15, 29, 4) {real, imag} */,
  {32'h4281fea0, 32'hc1b511fe} /* (15, 29, 3) {real, imag} */,
  {32'hc3e7a030, 32'hc2b40424} /* (15, 29, 2) {real, imag} */,
  {32'h44219be3, 32'h43c580ec} /* (15, 29, 1) {real, imag} */,
  {32'h448139eb, 32'h00000000} /* (15, 29, 0) {real, imag} */,
  {32'h43fb7a4e, 32'hc3b3ddfa} /* (15, 28, 31) {real, imag} */,
  {32'hc3f731fd, 32'hc2a57706} /* (15, 28, 30) {real, imag} */,
  {32'h426cd4b7, 32'h3e087400} /* (15, 28, 29) {real, imag} */,
  {32'h41abf5ee, 32'hc30f4b4e} /* (15, 28, 28) {real, imag} */,
  {32'hc2cb0493, 32'h422ec338} /* (15, 28, 27) {real, imag} */,
  {32'h42d27ad8, 32'h420ac7ca} /* (15, 28, 26) {real, imag} */,
  {32'h42fcd1cf, 32'hc2c9dd50} /* (15, 28, 25) {real, imag} */,
  {32'hc1ffbf3e, 32'hc153d634} /* (15, 28, 24) {real, imag} */,
  {32'h428f6232, 32'h4266a617} /* (15, 28, 23) {real, imag} */,
  {32'h4139e718, 32'hc00ead36} /* (15, 28, 22) {real, imag} */,
  {32'hc0456d2c, 32'hc108a324} /* (15, 28, 21) {real, imag} */,
  {32'h421bba95, 32'hc12a68f8} /* (15, 28, 20) {real, imag} */,
  {32'h41b1c2ec, 32'h42e51528} /* (15, 28, 19) {real, imag} */,
  {32'hc26a0bf8, 32'h423321cc} /* (15, 28, 18) {real, imag} */,
  {32'hc0ac8588, 32'hc1911792} /* (15, 28, 17) {real, imag} */,
  {32'h4206e4a5, 32'h00000000} /* (15, 28, 16) {real, imag} */,
  {32'hc0ac8588, 32'h41911792} /* (15, 28, 15) {real, imag} */,
  {32'hc26a0bf8, 32'hc23321cc} /* (15, 28, 14) {real, imag} */,
  {32'h41b1c2ec, 32'hc2e51528} /* (15, 28, 13) {real, imag} */,
  {32'h421bba95, 32'h412a68f8} /* (15, 28, 12) {real, imag} */,
  {32'hc0456d2c, 32'h4108a324} /* (15, 28, 11) {real, imag} */,
  {32'h4139e718, 32'h400ead36} /* (15, 28, 10) {real, imag} */,
  {32'h428f6232, 32'hc266a617} /* (15, 28, 9) {real, imag} */,
  {32'hc1ffbf3e, 32'h4153d634} /* (15, 28, 8) {real, imag} */,
  {32'h42fcd1cf, 32'h42c9dd50} /* (15, 28, 7) {real, imag} */,
  {32'h42d27ad8, 32'hc20ac7ca} /* (15, 28, 6) {real, imag} */,
  {32'hc2cb0493, 32'hc22ec338} /* (15, 28, 5) {real, imag} */,
  {32'h41abf5ee, 32'h430f4b4e} /* (15, 28, 4) {real, imag} */,
  {32'h426cd4b7, 32'hbe087400} /* (15, 28, 3) {real, imag} */,
  {32'hc3f731fd, 32'h42a57706} /* (15, 28, 2) {real, imag} */,
  {32'h43fb7a4e, 32'h43b3ddfa} /* (15, 28, 1) {real, imag} */,
  {32'h448c8bf4, 32'h00000000} /* (15, 28, 0) {real, imag} */,
  {32'h442b0ecd, 32'hc388243c} /* (15, 27, 31) {real, imag} */,
  {32'hc413b8b3, 32'hc1550fa8} /* (15, 27, 30) {real, imag} */,
  {32'h42d17999, 32'hc00a74e0} /* (15, 27, 29) {real, imag} */,
  {32'hc20cebda, 32'hc2f5ea5f} /* (15, 27, 28) {real, imag} */,
  {32'hbf0ebc00, 32'hc1b8e924} /* (15, 27, 27) {real, imag} */,
  {32'h42a6033d, 32'hc2b42f29} /* (15, 27, 26) {real, imag} */,
  {32'hc173e900, 32'hc22600ff} /* (15, 27, 25) {real, imag} */,
  {32'hc3105b01, 32'h43500dbc} /* (15, 27, 24) {real, imag} */,
  {32'h42a1081c, 32'hc1c10168} /* (15, 27, 23) {real, imag} */,
  {32'hc2983985, 32'hc274b499} /* (15, 27, 22) {real, imag} */,
  {32'hc18c6746, 32'h4127a234} /* (15, 27, 21) {real, imag} */,
  {32'h423a0b3f, 32'hc1e82b58} /* (15, 27, 20) {real, imag} */,
  {32'hc2229878, 32'h418ce1f4} /* (15, 27, 19) {real, imag} */,
  {32'h42a6cf78, 32'h42d9914d} /* (15, 27, 18) {real, imag} */,
  {32'hc032de70, 32'hc24c73a8} /* (15, 27, 17) {real, imag} */,
  {32'hc10cd290, 32'h00000000} /* (15, 27, 16) {real, imag} */,
  {32'hc032de70, 32'h424c73a8} /* (15, 27, 15) {real, imag} */,
  {32'h42a6cf78, 32'hc2d9914d} /* (15, 27, 14) {real, imag} */,
  {32'hc2229878, 32'hc18ce1f4} /* (15, 27, 13) {real, imag} */,
  {32'h423a0b3f, 32'h41e82b58} /* (15, 27, 12) {real, imag} */,
  {32'hc18c6746, 32'hc127a234} /* (15, 27, 11) {real, imag} */,
  {32'hc2983985, 32'h4274b499} /* (15, 27, 10) {real, imag} */,
  {32'h42a1081c, 32'h41c10168} /* (15, 27, 9) {real, imag} */,
  {32'hc3105b01, 32'hc3500dbc} /* (15, 27, 8) {real, imag} */,
  {32'hc173e900, 32'h422600ff} /* (15, 27, 7) {real, imag} */,
  {32'h42a6033d, 32'h42b42f29} /* (15, 27, 6) {real, imag} */,
  {32'hbf0ebc00, 32'h41b8e924} /* (15, 27, 5) {real, imag} */,
  {32'hc20cebda, 32'h42f5ea5f} /* (15, 27, 4) {real, imag} */,
  {32'h42d17999, 32'h400a74e0} /* (15, 27, 3) {real, imag} */,
  {32'hc413b8b3, 32'h41550fa8} /* (15, 27, 2) {real, imag} */,
  {32'h442b0ecd, 32'h4388243c} /* (15, 27, 1) {real, imag} */,
  {32'h446ee5d8, 32'h00000000} /* (15, 27, 0) {real, imag} */,
  {32'h445d5fe5, 32'hc338feec} /* (15, 26, 31) {real, imag} */,
  {32'hc401f138, 32'h41f121fc} /* (15, 26, 30) {real, imag} */,
  {32'h421e87b8, 32'h40198370} /* (15, 26, 29) {real, imag} */,
  {32'hc2f11124, 32'hc2e6279a} /* (15, 26, 28) {real, imag} */,
  {32'hc29385e7, 32'h433592d1} /* (15, 26, 27) {real, imag} */,
  {32'hc0be2c58, 32'hc28bb38c} /* (15, 26, 26) {real, imag} */,
  {32'hc1e06000, 32'h41e856f5} /* (15, 26, 25) {real, imag} */,
  {32'hc31aeb51, 32'hc1cbab42} /* (15, 26, 24) {real, imag} */,
  {32'h42af823f, 32'hc1a8415a} /* (15, 26, 23) {real, imag} */,
  {32'h429b233e, 32'hc2e601e8} /* (15, 26, 22) {real, imag} */,
  {32'h40d0cccc, 32'h42d00388} /* (15, 26, 21) {real, imag} */,
  {32'hc0e8ccd4, 32'hc2887d42} /* (15, 26, 20) {real, imag} */,
  {32'h42095504, 32'h4192903a} /* (15, 26, 19) {real, imag} */,
  {32'h42b9dbc0, 32'h42816d5f} /* (15, 26, 18) {real, imag} */,
  {32'h420039c6, 32'hc1c97be6} /* (15, 26, 17) {real, imag} */,
  {32'hc1d45a26, 32'h00000000} /* (15, 26, 16) {real, imag} */,
  {32'h420039c6, 32'h41c97be6} /* (15, 26, 15) {real, imag} */,
  {32'h42b9dbc0, 32'hc2816d5f} /* (15, 26, 14) {real, imag} */,
  {32'h42095504, 32'hc192903a} /* (15, 26, 13) {real, imag} */,
  {32'hc0e8ccd4, 32'h42887d42} /* (15, 26, 12) {real, imag} */,
  {32'h40d0cccc, 32'hc2d00388} /* (15, 26, 11) {real, imag} */,
  {32'h429b233e, 32'h42e601e8} /* (15, 26, 10) {real, imag} */,
  {32'h42af823f, 32'h41a8415a} /* (15, 26, 9) {real, imag} */,
  {32'hc31aeb51, 32'h41cbab42} /* (15, 26, 8) {real, imag} */,
  {32'hc1e06000, 32'hc1e856f5} /* (15, 26, 7) {real, imag} */,
  {32'hc0be2c58, 32'h428bb38c} /* (15, 26, 6) {real, imag} */,
  {32'hc29385e7, 32'hc33592d1} /* (15, 26, 5) {real, imag} */,
  {32'hc2f11124, 32'h42e6279a} /* (15, 26, 4) {real, imag} */,
  {32'h421e87b8, 32'hc0198370} /* (15, 26, 3) {real, imag} */,
  {32'hc401f138, 32'hc1f121fc} /* (15, 26, 2) {real, imag} */,
  {32'h445d5fe5, 32'h4338feec} /* (15, 26, 1) {real, imag} */,
  {32'h443204a4, 32'h00000000} /* (15, 26, 0) {real, imag} */,
  {32'h44673852, 32'hc31b54ae} /* (15, 25, 31) {real, imag} */,
  {32'hc401c6d3, 32'h42d34958} /* (15, 25, 30) {real, imag} */,
  {32'h42a23f34, 32'hc2ae5d63} /* (15, 25, 29) {real, imag} */,
  {32'h40c8b8d8, 32'hc1f722f4} /* (15, 25, 28) {real, imag} */,
  {32'hc272da65, 32'h430a163e} /* (15, 25, 27) {real, imag} */,
  {32'h42a90978, 32'h41c43edb} /* (15, 25, 26) {real, imag} */,
  {32'h421e3894, 32'h426e4250} /* (15, 25, 25) {real, imag} */,
  {32'hc0bf1c14, 32'h41244ba4} /* (15, 25, 24) {real, imag} */,
  {32'h42a5253a, 32'h42688a4e} /* (15, 25, 23) {real, imag} */,
  {32'hc23eac7c, 32'h42940fe2} /* (15, 25, 22) {real, imag} */,
  {32'h41c1a147, 32'hc220e0f0} /* (15, 25, 21) {real, imag} */,
  {32'hc1046faa, 32'h4249e11b} /* (15, 25, 20) {real, imag} */,
  {32'hc22b9808, 32'h41192d48} /* (15, 25, 19) {real, imag} */,
  {32'hc262412a, 32'h42805ecd} /* (15, 25, 18) {real, imag} */,
  {32'hc14c269f, 32'hc1a2dc87} /* (15, 25, 17) {real, imag} */,
  {32'hbf4a1d20, 32'h00000000} /* (15, 25, 16) {real, imag} */,
  {32'hc14c269f, 32'h41a2dc87} /* (15, 25, 15) {real, imag} */,
  {32'hc262412a, 32'hc2805ecd} /* (15, 25, 14) {real, imag} */,
  {32'hc22b9808, 32'hc1192d48} /* (15, 25, 13) {real, imag} */,
  {32'hc1046faa, 32'hc249e11b} /* (15, 25, 12) {real, imag} */,
  {32'h41c1a147, 32'h4220e0f0} /* (15, 25, 11) {real, imag} */,
  {32'hc23eac7c, 32'hc2940fe2} /* (15, 25, 10) {real, imag} */,
  {32'h42a5253a, 32'hc2688a4e} /* (15, 25, 9) {real, imag} */,
  {32'hc0bf1c14, 32'hc1244ba4} /* (15, 25, 8) {real, imag} */,
  {32'h421e3894, 32'hc26e4250} /* (15, 25, 7) {real, imag} */,
  {32'h42a90978, 32'hc1c43edb} /* (15, 25, 6) {real, imag} */,
  {32'hc272da65, 32'hc30a163e} /* (15, 25, 5) {real, imag} */,
  {32'h40c8b8d8, 32'h41f722f4} /* (15, 25, 4) {real, imag} */,
  {32'h42a23f34, 32'h42ae5d63} /* (15, 25, 3) {real, imag} */,
  {32'hc401c6d3, 32'hc2d34958} /* (15, 25, 2) {real, imag} */,
  {32'h44673852, 32'h431b54ae} /* (15, 25, 1) {real, imag} */,
  {32'h4433a4de, 32'h00000000} /* (15, 25, 0) {real, imag} */,
  {32'h44592fe9, 32'hc343af4f} /* (15, 24, 31) {real, imag} */,
  {32'hc3dce43d, 32'h43103cb2} /* (15, 24, 30) {real, imag} */,
  {32'h428c1ced, 32'hc31e20ce} /* (15, 24, 29) {real, imag} */,
  {32'h4073dfa8, 32'hc3135650} /* (15, 24, 28) {real, imag} */,
  {32'hc2b9b116, 32'h41da2f94} /* (15, 24, 27) {real, imag} */,
  {32'hc29ed456, 32'h43118c05} /* (15, 24, 26) {real, imag} */,
  {32'h429103cc, 32'hc1fd96bc} /* (15, 24, 25) {real, imag} */,
  {32'h4215d722, 32'h424de0dd} /* (15, 24, 24) {real, imag} */,
  {32'hc28571fa, 32'hc118eb8c} /* (15, 24, 23) {real, imag} */,
  {32'hc0e34d78, 32'hc261776e} /* (15, 24, 22) {real, imag} */,
  {32'h4230716b, 32'h4277e8da} /* (15, 24, 21) {real, imag} */,
  {32'hc24bf9d9, 32'hc15e2040} /* (15, 24, 20) {real, imag} */,
  {32'h4242669e, 32'h41e7eecc} /* (15, 24, 19) {real, imag} */,
  {32'hc1b8fd05, 32'h423be2d0} /* (15, 24, 18) {real, imag} */,
  {32'hc182ef72, 32'hc1dd99ad} /* (15, 24, 17) {real, imag} */,
  {32'h4261ad94, 32'h00000000} /* (15, 24, 16) {real, imag} */,
  {32'hc182ef72, 32'h41dd99ad} /* (15, 24, 15) {real, imag} */,
  {32'hc1b8fd05, 32'hc23be2d0} /* (15, 24, 14) {real, imag} */,
  {32'h4242669e, 32'hc1e7eecc} /* (15, 24, 13) {real, imag} */,
  {32'hc24bf9d9, 32'h415e2040} /* (15, 24, 12) {real, imag} */,
  {32'h4230716b, 32'hc277e8da} /* (15, 24, 11) {real, imag} */,
  {32'hc0e34d78, 32'h4261776e} /* (15, 24, 10) {real, imag} */,
  {32'hc28571fa, 32'h4118eb8c} /* (15, 24, 9) {real, imag} */,
  {32'h4215d722, 32'hc24de0dd} /* (15, 24, 8) {real, imag} */,
  {32'h429103cc, 32'h41fd96bc} /* (15, 24, 7) {real, imag} */,
  {32'hc29ed456, 32'hc3118c05} /* (15, 24, 6) {real, imag} */,
  {32'hc2b9b116, 32'hc1da2f94} /* (15, 24, 5) {real, imag} */,
  {32'h4073dfa8, 32'h43135650} /* (15, 24, 4) {real, imag} */,
  {32'h428c1ced, 32'h431e20ce} /* (15, 24, 3) {real, imag} */,
  {32'hc3dce43d, 32'hc3103cb2} /* (15, 24, 2) {real, imag} */,
  {32'h44592fe9, 32'h4343af4f} /* (15, 24, 1) {real, imag} */,
  {32'h4410f00c, 32'h00000000} /* (15, 24, 0) {real, imag} */,
  {32'h44431bac, 32'hc2cdeec1} /* (15, 23, 31) {real, imag} */,
  {32'hc3cdfb6a, 32'h42e7a984} /* (15, 23, 30) {real, imag} */,
  {32'hc27b7788, 32'hc37ff318} /* (15, 23, 29) {real, imag} */,
  {32'hc2a625d8, 32'hc37f923a} /* (15, 23, 28) {real, imag} */,
  {32'hc3075132, 32'hc104575e} /* (15, 23, 27) {real, imag} */,
  {32'hc2e5f91c, 32'hc295428b} /* (15, 23, 26) {real, imag} */,
  {32'h4292ac85, 32'h421cf9b6} /* (15, 23, 25) {real, imag} */,
  {32'hc2128cc2, 32'h42c4c0f0} /* (15, 23, 24) {real, imag} */,
  {32'h424fbac5, 32'h408d384d} /* (15, 23, 23) {real, imag} */,
  {32'hc1ad8ec8, 32'h42388505} /* (15, 23, 22) {real, imag} */,
  {32'h408abc28, 32'h41af2405} /* (15, 23, 21) {real, imag} */,
  {32'h42002238, 32'hc2ad5abd} /* (15, 23, 20) {real, imag} */,
  {32'h3f9649a0, 32'hc288e62f} /* (15, 23, 19) {real, imag} */,
  {32'h42806b38, 32'h41c7db25} /* (15, 23, 18) {real, imag} */,
  {32'hc1bf50ea, 32'h42ba8019} /* (15, 23, 17) {real, imag} */,
  {32'hc3027801, 32'h00000000} /* (15, 23, 16) {real, imag} */,
  {32'hc1bf50ea, 32'hc2ba8019} /* (15, 23, 15) {real, imag} */,
  {32'h42806b38, 32'hc1c7db25} /* (15, 23, 14) {real, imag} */,
  {32'h3f9649a0, 32'h4288e62f} /* (15, 23, 13) {real, imag} */,
  {32'h42002238, 32'h42ad5abd} /* (15, 23, 12) {real, imag} */,
  {32'h408abc28, 32'hc1af2405} /* (15, 23, 11) {real, imag} */,
  {32'hc1ad8ec8, 32'hc2388505} /* (15, 23, 10) {real, imag} */,
  {32'h424fbac5, 32'hc08d384d} /* (15, 23, 9) {real, imag} */,
  {32'hc2128cc2, 32'hc2c4c0f0} /* (15, 23, 8) {real, imag} */,
  {32'h4292ac85, 32'hc21cf9b6} /* (15, 23, 7) {real, imag} */,
  {32'hc2e5f91c, 32'h4295428b} /* (15, 23, 6) {real, imag} */,
  {32'hc3075132, 32'h4104575e} /* (15, 23, 5) {real, imag} */,
  {32'hc2a625d8, 32'h437f923a} /* (15, 23, 4) {real, imag} */,
  {32'hc27b7788, 32'h437ff318} /* (15, 23, 3) {real, imag} */,
  {32'hc3cdfb6a, 32'hc2e7a984} /* (15, 23, 2) {real, imag} */,
  {32'h44431bac, 32'h42cdeec1} /* (15, 23, 1) {real, imag} */,
  {32'h43b0aa4d, 32'h00000000} /* (15, 23, 0) {real, imag} */,
  {32'h4428c32a, 32'hc2925339} /* (15, 22, 31) {real, imag} */,
  {32'hc381815a, 32'h42cec0c2} /* (15, 22, 30) {real, imag} */,
  {32'h424029de, 32'hc346ccb4} /* (15, 22, 29) {real, imag} */,
  {32'hc25925eb, 32'hc33db051} /* (15, 22, 28) {real, imag} */,
  {32'hc295f181, 32'h41928705} /* (15, 22, 27) {real, imag} */,
  {32'hc326517e, 32'hc296ea08} /* (15, 22, 26) {real, imag} */,
  {32'h42f16736, 32'h417e5e08} /* (15, 22, 25) {real, imag} */,
  {32'hc0ef4e40, 32'h420c27ba} /* (15, 22, 24) {real, imag} */,
  {32'hc12ca4ee, 32'h3f0e7570} /* (15, 22, 23) {real, imag} */,
  {32'hc2ddb5fe, 32'hc12fed48} /* (15, 22, 22) {real, imag} */,
  {32'hc20bb33f, 32'hc2051386} /* (15, 22, 21) {real, imag} */,
  {32'hc245d0de, 32'hc24a28ba} /* (15, 22, 20) {real, imag} */,
  {32'h40a02c20, 32'h41fd3214} /* (15, 22, 19) {real, imag} */,
  {32'hc29d165b, 32'h402be7b4} /* (15, 22, 18) {real, imag} */,
  {32'hbf645e80, 32'hc23672fb} /* (15, 22, 17) {real, imag} */,
  {32'h425aa288, 32'h00000000} /* (15, 22, 16) {real, imag} */,
  {32'hbf645e80, 32'h423672fb} /* (15, 22, 15) {real, imag} */,
  {32'hc29d165b, 32'hc02be7b4} /* (15, 22, 14) {real, imag} */,
  {32'h40a02c20, 32'hc1fd3214} /* (15, 22, 13) {real, imag} */,
  {32'hc245d0de, 32'h424a28ba} /* (15, 22, 12) {real, imag} */,
  {32'hc20bb33f, 32'h42051386} /* (15, 22, 11) {real, imag} */,
  {32'hc2ddb5fe, 32'h412fed48} /* (15, 22, 10) {real, imag} */,
  {32'hc12ca4ee, 32'hbf0e7570} /* (15, 22, 9) {real, imag} */,
  {32'hc0ef4e40, 32'hc20c27ba} /* (15, 22, 8) {real, imag} */,
  {32'h42f16736, 32'hc17e5e08} /* (15, 22, 7) {real, imag} */,
  {32'hc326517e, 32'h4296ea08} /* (15, 22, 6) {real, imag} */,
  {32'hc295f181, 32'hc1928705} /* (15, 22, 5) {real, imag} */,
  {32'hc25925eb, 32'h433db051} /* (15, 22, 4) {real, imag} */,
  {32'h424029de, 32'h4346ccb4} /* (15, 22, 3) {real, imag} */,
  {32'hc381815a, 32'hc2cec0c2} /* (15, 22, 2) {real, imag} */,
  {32'h4428c32a, 32'h42925339} /* (15, 22, 1) {real, imag} */,
  {32'h4372ccf4, 32'h00000000} /* (15, 22, 0) {real, imag} */,
  {32'h4341400a, 32'hc283f426} /* (15, 21, 31) {real, imag} */,
  {32'hc2a0ee8c, 32'h4301c91c} /* (15, 21, 30) {real, imag} */,
  {32'h428338b0, 32'hc2e8fede} /* (15, 21, 29) {real, imag} */,
  {32'h4198d1a0, 32'hc327a81b} /* (15, 21, 28) {real, imag} */,
  {32'hc2a0159b, 32'hc1139c40} /* (15, 21, 27) {real, imag} */,
  {32'h421a29d8, 32'hc20532a4} /* (15, 21, 26) {real, imag} */,
  {32'h4274e7e8, 32'h4146572c} /* (15, 21, 25) {real, imag} */,
  {32'hc24c2998, 32'hc21fd2e4} /* (15, 21, 24) {real, imag} */,
  {32'h418de962, 32'hc1c4289e} /* (15, 21, 23) {real, imag} */,
  {32'h414b04e8, 32'h4120c264} /* (15, 21, 22) {real, imag} */,
  {32'h420306c3, 32'h4308d8ff} /* (15, 21, 21) {real, imag} */,
  {32'hc14e3c18, 32'h42991cd5} /* (15, 21, 20) {real, imag} */,
  {32'h3fd190c0, 32'hc15579c4} /* (15, 21, 19) {real, imag} */,
  {32'hc0e1fdd2, 32'h4157d9b4} /* (15, 21, 18) {real, imag} */,
  {32'h42ad825e, 32'h41d3738a} /* (15, 21, 17) {real, imag} */,
  {32'hc14b8c78, 32'h00000000} /* (15, 21, 16) {real, imag} */,
  {32'h42ad825e, 32'hc1d3738a} /* (15, 21, 15) {real, imag} */,
  {32'hc0e1fdd2, 32'hc157d9b4} /* (15, 21, 14) {real, imag} */,
  {32'h3fd190c0, 32'h415579c4} /* (15, 21, 13) {real, imag} */,
  {32'hc14e3c18, 32'hc2991cd5} /* (15, 21, 12) {real, imag} */,
  {32'h420306c3, 32'hc308d8ff} /* (15, 21, 11) {real, imag} */,
  {32'h414b04e8, 32'hc120c264} /* (15, 21, 10) {real, imag} */,
  {32'h418de962, 32'h41c4289e} /* (15, 21, 9) {real, imag} */,
  {32'hc24c2998, 32'h421fd2e4} /* (15, 21, 8) {real, imag} */,
  {32'h4274e7e8, 32'hc146572c} /* (15, 21, 7) {real, imag} */,
  {32'h421a29d8, 32'h420532a4} /* (15, 21, 6) {real, imag} */,
  {32'hc2a0159b, 32'h41139c40} /* (15, 21, 5) {real, imag} */,
  {32'h4198d1a0, 32'h4327a81b} /* (15, 21, 4) {real, imag} */,
  {32'h428338b0, 32'h42e8fede} /* (15, 21, 3) {real, imag} */,
  {32'hc2a0ee8c, 32'hc301c91c} /* (15, 21, 2) {real, imag} */,
  {32'h4341400a, 32'h4283f426} /* (15, 21, 1) {real, imag} */,
  {32'hc1190d70, 32'h00000000} /* (15, 21, 0) {real, imag} */,
  {32'hc3fe2f3a, 32'h433d83b2} /* (15, 20, 31) {real, imag} */,
  {32'h4386ae06, 32'hc0705eb0} /* (15, 20, 30) {real, imag} */,
  {32'h43077f14, 32'hc1831678} /* (15, 20, 29) {real, imag} */,
  {32'h407a8b00, 32'hc27edd4a} /* (15, 20, 28) {real, imag} */,
  {32'h41cf1f03, 32'h3f512f80} /* (15, 20, 27) {real, imag} */,
  {32'hc178af2c, 32'hc29325ca} /* (15, 20, 26) {real, imag} */,
  {32'hc30c6aa2, 32'hc22d2df5} /* (15, 20, 25) {real, imag} */,
  {32'h42b05210, 32'hc305a20f} /* (15, 20, 24) {real, imag} */,
  {32'h41db45c2, 32'h420c7d26} /* (15, 20, 23) {real, imag} */,
  {32'h41802615, 32'hc14626c4} /* (15, 20, 22) {real, imag} */,
  {32'hc2108b43, 32'hc1d13ca0} /* (15, 20, 21) {real, imag} */,
  {32'hc25a6054, 32'h42072aba} /* (15, 20, 20) {real, imag} */,
  {32'hc21b196a, 32'hc250e24d} /* (15, 20, 19) {real, imag} */,
  {32'hc12fc2b2, 32'hc1d29695} /* (15, 20, 18) {real, imag} */,
  {32'h412c5c15, 32'hbff10470} /* (15, 20, 17) {real, imag} */,
  {32'h41d41e39, 32'h00000000} /* (15, 20, 16) {real, imag} */,
  {32'h412c5c15, 32'h3ff10470} /* (15, 20, 15) {real, imag} */,
  {32'hc12fc2b2, 32'h41d29695} /* (15, 20, 14) {real, imag} */,
  {32'hc21b196a, 32'h4250e24d} /* (15, 20, 13) {real, imag} */,
  {32'hc25a6054, 32'hc2072aba} /* (15, 20, 12) {real, imag} */,
  {32'hc2108b43, 32'h41d13ca0} /* (15, 20, 11) {real, imag} */,
  {32'h41802615, 32'h414626c4} /* (15, 20, 10) {real, imag} */,
  {32'h41db45c2, 32'hc20c7d26} /* (15, 20, 9) {real, imag} */,
  {32'h42b05210, 32'h4305a20f} /* (15, 20, 8) {real, imag} */,
  {32'hc30c6aa2, 32'h422d2df5} /* (15, 20, 7) {real, imag} */,
  {32'hc178af2c, 32'h429325ca} /* (15, 20, 6) {real, imag} */,
  {32'h41cf1f03, 32'hbf512f80} /* (15, 20, 5) {real, imag} */,
  {32'h407a8b00, 32'h427edd4a} /* (15, 20, 4) {real, imag} */,
  {32'h43077f14, 32'h41831678} /* (15, 20, 3) {real, imag} */,
  {32'h4386ae06, 32'h40705eb0} /* (15, 20, 2) {real, imag} */,
  {32'hc3fe2f3a, 32'hc33d83b2} /* (15, 20, 1) {real, imag} */,
  {32'hc3af4937, 32'h00000000} /* (15, 20, 0) {real, imag} */,
  {32'hc446a411, 32'h4356fe53} /* (15, 19, 31) {real, imag} */,
  {32'h43c305e4, 32'hc224f326} /* (15, 19, 30) {real, imag} */,
  {32'h4323f84c, 32'h42132e34} /* (15, 19, 29) {real, imag} */,
  {32'h420aa5ca, 32'hc2ee9eb8} /* (15, 19, 28) {real, imag} */,
  {32'h429bbe62, 32'h42077249} /* (15, 19, 27) {real, imag} */,
  {32'hc2b251c2, 32'hc18299ce} /* (15, 19, 26) {real, imag} */,
  {32'hc2b49dac, 32'h41dacf6a} /* (15, 19, 25) {real, imag} */,
  {32'h42107490, 32'hc21441e5} /* (15, 19, 24) {real, imag} */,
  {32'hc2e7a634, 32'h4101d840} /* (15, 19, 23) {real, imag} */,
  {32'h40f10770, 32'hc28cba73} /* (15, 19, 22) {real, imag} */,
  {32'h41236f72, 32'hc2ac8390} /* (15, 19, 21) {real, imag} */,
  {32'h42793aa1, 32'hc29311da} /* (15, 19, 20) {real, imag} */,
  {32'hc1aab737, 32'h41e30b34} /* (15, 19, 19) {real, imag} */,
  {32'hc18a9b26, 32'h42b534fc} /* (15, 19, 18) {real, imag} */,
  {32'h4147f7b4, 32'h42871996} /* (15, 19, 17) {real, imag} */,
  {32'hc07bc984, 32'h00000000} /* (15, 19, 16) {real, imag} */,
  {32'h4147f7b4, 32'hc2871996} /* (15, 19, 15) {real, imag} */,
  {32'hc18a9b26, 32'hc2b534fc} /* (15, 19, 14) {real, imag} */,
  {32'hc1aab737, 32'hc1e30b34} /* (15, 19, 13) {real, imag} */,
  {32'h42793aa1, 32'h429311da} /* (15, 19, 12) {real, imag} */,
  {32'h41236f72, 32'h42ac8390} /* (15, 19, 11) {real, imag} */,
  {32'h40f10770, 32'h428cba73} /* (15, 19, 10) {real, imag} */,
  {32'hc2e7a634, 32'hc101d840} /* (15, 19, 9) {real, imag} */,
  {32'h42107490, 32'h421441e5} /* (15, 19, 8) {real, imag} */,
  {32'hc2b49dac, 32'hc1dacf6a} /* (15, 19, 7) {real, imag} */,
  {32'hc2b251c2, 32'h418299ce} /* (15, 19, 6) {real, imag} */,
  {32'h429bbe62, 32'hc2077249} /* (15, 19, 5) {real, imag} */,
  {32'h420aa5ca, 32'h42ee9eb8} /* (15, 19, 4) {real, imag} */,
  {32'h4323f84c, 32'hc2132e34} /* (15, 19, 3) {real, imag} */,
  {32'h43c305e4, 32'h4224f326} /* (15, 19, 2) {real, imag} */,
  {32'hc446a411, 32'hc356fe53} /* (15, 19, 1) {real, imag} */,
  {32'hc3c64828, 32'h00000000} /* (15, 19, 0) {real, imag} */,
  {32'hc454672b, 32'h422481a8} /* (15, 18, 31) {real, imag} */,
  {32'h43d0d966, 32'hc210af02} /* (15, 18, 30) {real, imag} */,
  {32'h430f1c6e, 32'h42981aae} /* (15, 18, 29) {real, imag} */,
  {32'hc3055fb3, 32'h4338c1e2} /* (15, 18, 28) {real, imag} */,
  {32'h42aee1ba, 32'hc30d160f} /* (15, 18, 27) {real, imag} */,
  {32'hc1ff0174, 32'hc20a85fa} /* (15, 18, 26) {real, imag} */,
  {32'h415db750, 32'hc1c2c01a} /* (15, 18, 25) {real, imag} */,
  {32'h42d11bfd, 32'h42b5aa63} /* (15, 18, 24) {real, imag} */,
  {32'h418ca675, 32'hc13ef9ce} /* (15, 18, 23) {real, imag} */,
  {32'hc2c69bf1, 32'h41b60afc} /* (15, 18, 22) {real, imag} */,
  {32'hc0920bb4, 32'h42b38f5a} /* (15, 18, 21) {real, imag} */,
  {32'h425774fc, 32'hc2385dce} /* (15, 18, 20) {real, imag} */,
  {32'hc29e4911, 32'hc201a46c} /* (15, 18, 19) {real, imag} */,
  {32'hc27b66f9, 32'hc26b3cb4} /* (15, 18, 18) {real, imag} */,
  {32'hc1e38901, 32'hc18612db} /* (15, 18, 17) {real, imag} */,
  {32'hc1b1e30f, 32'h00000000} /* (15, 18, 16) {real, imag} */,
  {32'hc1e38901, 32'h418612db} /* (15, 18, 15) {real, imag} */,
  {32'hc27b66f9, 32'h426b3cb4} /* (15, 18, 14) {real, imag} */,
  {32'hc29e4911, 32'h4201a46c} /* (15, 18, 13) {real, imag} */,
  {32'h425774fc, 32'h42385dce} /* (15, 18, 12) {real, imag} */,
  {32'hc0920bb4, 32'hc2b38f5a} /* (15, 18, 11) {real, imag} */,
  {32'hc2c69bf1, 32'hc1b60afc} /* (15, 18, 10) {real, imag} */,
  {32'h418ca675, 32'h413ef9ce} /* (15, 18, 9) {real, imag} */,
  {32'h42d11bfd, 32'hc2b5aa63} /* (15, 18, 8) {real, imag} */,
  {32'h415db750, 32'h41c2c01a} /* (15, 18, 7) {real, imag} */,
  {32'hc1ff0174, 32'h420a85fa} /* (15, 18, 6) {real, imag} */,
  {32'h42aee1ba, 32'h430d160f} /* (15, 18, 5) {real, imag} */,
  {32'hc3055fb3, 32'hc338c1e2} /* (15, 18, 4) {real, imag} */,
  {32'h430f1c6e, 32'hc2981aae} /* (15, 18, 3) {real, imag} */,
  {32'h43d0d966, 32'h4210af02} /* (15, 18, 2) {real, imag} */,
  {32'hc454672b, 32'hc22481a8} /* (15, 18, 1) {real, imag} */,
  {32'hc3f5b7dc, 32'h00000000} /* (15, 18, 0) {real, imag} */,
  {32'hc46a0e51, 32'h42053c50} /* (15, 17, 31) {real, imag} */,
  {32'h43f270dd, 32'hbff31620} /* (15, 17, 30) {real, imag} */,
  {32'h42b9067e, 32'hc207b67a} /* (15, 17, 29) {real, imag} */,
  {32'hc1c936fe, 32'h43363b93} /* (15, 17, 28) {real, imag} */,
  {32'h418be5be, 32'hc294f4ba} /* (15, 17, 27) {real, imag} */,
  {32'hc2d8ef95, 32'h4281df82} /* (15, 17, 26) {real, imag} */,
  {32'hc2db05d0, 32'hc20bd1b3} /* (15, 17, 25) {real, imag} */,
  {32'h4307a58b, 32'hc294abe8} /* (15, 17, 24) {real, imag} */,
  {32'h418065bc, 32'h415268a2} /* (15, 17, 23) {real, imag} */,
  {32'hc2b6a4c8, 32'hc139ba76} /* (15, 17, 22) {real, imag} */,
  {32'h42258172, 32'hc274ce8e} /* (15, 17, 21) {real, imag} */,
  {32'hc286d39e, 32'hc2867952} /* (15, 17, 20) {real, imag} */,
  {32'hc19f4e52, 32'hc2103a6e} /* (15, 17, 19) {real, imag} */,
  {32'hc16cdfd4, 32'h416db26c} /* (15, 17, 18) {real, imag} */,
  {32'h40915aa8, 32'h4204245d} /* (15, 17, 17) {real, imag} */,
  {32'hc24b82c8, 32'h00000000} /* (15, 17, 16) {real, imag} */,
  {32'h40915aa8, 32'hc204245d} /* (15, 17, 15) {real, imag} */,
  {32'hc16cdfd4, 32'hc16db26c} /* (15, 17, 14) {real, imag} */,
  {32'hc19f4e52, 32'h42103a6e} /* (15, 17, 13) {real, imag} */,
  {32'hc286d39e, 32'h42867952} /* (15, 17, 12) {real, imag} */,
  {32'h42258172, 32'h4274ce8e} /* (15, 17, 11) {real, imag} */,
  {32'hc2b6a4c8, 32'h4139ba76} /* (15, 17, 10) {real, imag} */,
  {32'h418065bc, 32'hc15268a2} /* (15, 17, 9) {real, imag} */,
  {32'h4307a58b, 32'h4294abe8} /* (15, 17, 8) {real, imag} */,
  {32'hc2db05d0, 32'h420bd1b3} /* (15, 17, 7) {real, imag} */,
  {32'hc2d8ef95, 32'hc281df82} /* (15, 17, 6) {real, imag} */,
  {32'h418be5be, 32'h4294f4ba} /* (15, 17, 5) {real, imag} */,
  {32'hc1c936fe, 32'hc3363b93} /* (15, 17, 4) {real, imag} */,
  {32'h42b9067e, 32'h4207b67a} /* (15, 17, 3) {real, imag} */,
  {32'h43f270dd, 32'h3ff31620} /* (15, 17, 2) {real, imag} */,
  {32'hc46a0e51, 32'hc2053c50} /* (15, 17, 1) {real, imag} */,
  {32'hc4439a26, 32'h00000000} /* (15, 17, 0) {real, imag} */,
  {32'hc4801cb5, 32'h434e78f5} /* (15, 16, 31) {real, imag} */,
  {32'h440b1472, 32'h4101f5c0} /* (15, 16, 30) {real, imag} */,
  {32'h434658f0, 32'hc2dd41af} /* (15, 16, 29) {real, imag} */,
  {32'hc31134f6, 32'h434cb82d} /* (15, 16, 28) {real, imag} */,
  {32'hc16be700, 32'hc28e0496} /* (15, 16, 27) {real, imag} */,
  {32'hc2ba2096, 32'h41427c90} /* (15, 16, 26) {real, imag} */,
  {32'h42cced87, 32'h4150d0b5} /* (15, 16, 25) {real, imag} */,
  {32'h4293cbcc, 32'hc20caf2b} /* (15, 16, 24) {real, imag} */,
  {32'h423b2579, 32'hc24da6a5} /* (15, 16, 23) {real, imag} */,
  {32'h41bc2deb, 32'hc123f363} /* (15, 16, 22) {real, imag} */,
  {32'h42281104, 32'hc229ede4} /* (15, 16, 21) {real, imag} */,
  {32'hc22e6dba, 32'hc2630a9d} /* (15, 16, 20) {real, imag} */,
  {32'hc21739f3, 32'h423f56b3} /* (15, 16, 19) {real, imag} */,
  {32'h41b6b077, 32'h420d5739} /* (15, 16, 18) {real, imag} */,
  {32'h421839c4, 32'hc130370e} /* (15, 16, 17) {real, imag} */,
  {32'h413201ca, 32'h00000000} /* (15, 16, 16) {real, imag} */,
  {32'h421839c4, 32'h4130370e} /* (15, 16, 15) {real, imag} */,
  {32'h41b6b077, 32'hc20d5739} /* (15, 16, 14) {real, imag} */,
  {32'hc21739f3, 32'hc23f56b3} /* (15, 16, 13) {real, imag} */,
  {32'hc22e6dba, 32'h42630a9d} /* (15, 16, 12) {real, imag} */,
  {32'h42281104, 32'h4229ede4} /* (15, 16, 11) {real, imag} */,
  {32'h41bc2deb, 32'h4123f363} /* (15, 16, 10) {real, imag} */,
  {32'h423b2579, 32'h424da6a5} /* (15, 16, 9) {real, imag} */,
  {32'h4293cbcc, 32'h420caf2b} /* (15, 16, 8) {real, imag} */,
  {32'h42cced87, 32'hc150d0b5} /* (15, 16, 7) {real, imag} */,
  {32'hc2ba2096, 32'hc1427c90} /* (15, 16, 6) {real, imag} */,
  {32'hc16be700, 32'h428e0496} /* (15, 16, 5) {real, imag} */,
  {32'hc31134f6, 32'hc34cb82d} /* (15, 16, 4) {real, imag} */,
  {32'h434658f0, 32'h42dd41af} /* (15, 16, 3) {real, imag} */,
  {32'h440b1472, 32'hc101f5c0} /* (15, 16, 2) {real, imag} */,
  {32'hc4801cb5, 32'hc34e78f5} /* (15, 16, 1) {real, imag} */,
  {32'hc458b48d, 32'h00000000} /* (15, 16, 0) {real, imag} */,
  {32'hc493541e, 32'h4386a81a} /* (15, 15, 31) {real, imag} */,
  {32'h440f65ad, 32'h4096bae8} /* (15, 15, 30) {real, imag} */,
  {32'h4303d352, 32'hc2c7d28f} /* (15, 15, 29) {real, imag} */,
  {32'hc300caf7, 32'h42b2c5aa} /* (15, 15, 28) {real, imag} */,
  {32'hc2664d59, 32'hc2248938} /* (15, 15, 27) {real, imag} */,
  {32'hc2696dee, 32'h43011453} /* (15, 15, 26) {real, imag} */,
  {32'h420c1d0c, 32'hc209f29d} /* (15, 15, 25) {real, imag} */,
  {32'h4285951e, 32'hc21fea6d} /* (15, 15, 24) {real, imag} */,
  {32'h42983181, 32'hc1d03659} /* (15, 15, 23) {real, imag} */,
  {32'hc1894f30, 32'h408ea6ec} /* (15, 15, 22) {real, imag} */,
  {32'hc02e0a18, 32'h425114a6} /* (15, 15, 21) {real, imag} */,
  {32'h42ae2112, 32'hc2769e44} /* (15, 15, 20) {real, imag} */,
  {32'hc2d9982a, 32'h422b70a8} /* (15, 15, 19) {real, imag} */,
  {32'h425e7269, 32'hc1c36260} /* (15, 15, 18) {real, imag} */,
  {32'hc211d0c1, 32'hc20da55b} /* (15, 15, 17) {real, imag} */,
  {32'h4145b216, 32'h00000000} /* (15, 15, 16) {real, imag} */,
  {32'hc211d0c1, 32'h420da55b} /* (15, 15, 15) {real, imag} */,
  {32'h425e7269, 32'h41c36260} /* (15, 15, 14) {real, imag} */,
  {32'hc2d9982a, 32'hc22b70a8} /* (15, 15, 13) {real, imag} */,
  {32'h42ae2112, 32'h42769e44} /* (15, 15, 12) {real, imag} */,
  {32'hc02e0a18, 32'hc25114a6} /* (15, 15, 11) {real, imag} */,
  {32'hc1894f30, 32'hc08ea6ec} /* (15, 15, 10) {real, imag} */,
  {32'h42983181, 32'h41d03659} /* (15, 15, 9) {real, imag} */,
  {32'h4285951e, 32'h421fea6d} /* (15, 15, 8) {real, imag} */,
  {32'h420c1d0c, 32'h4209f29d} /* (15, 15, 7) {real, imag} */,
  {32'hc2696dee, 32'hc3011453} /* (15, 15, 6) {real, imag} */,
  {32'hc2664d59, 32'h42248938} /* (15, 15, 5) {real, imag} */,
  {32'hc300caf7, 32'hc2b2c5aa} /* (15, 15, 4) {real, imag} */,
  {32'h4303d352, 32'h42c7d28f} /* (15, 15, 3) {real, imag} */,
  {32'h440f65ad, 32'hc096bae8} /* (15, 15, 2) {real, imag} */,
  {32'hc493541e, 32'hc386a81a} /* (15, 15, 1) {real, imag} */,
  {32'hc431085a, 32'h00000000} /* (15, 15, 0) {real, imag} */,
  {32'hc4a31fed, 32'h43e1bec1} /* (15, 14, 31) {real, imag} */,
  {32'h44023bfd, 32'h42b83523} /* (15, 14, 30) {real, imag} */,
  {32'h43274f4e, 32'hc18a35fa} /* (15, 14, 29) {real, imag} */,
  {32'hc217590c, 32'h4321be90} /* (15, 14, 28) {real, imag} */,
  {32'h4035dc90, 32'hc3128fed} /* (15, 14, 27) {real, imag} */,
  {32'h41b8cdc8, 32'hc2188bc8} /* (15, 14, 26) {real, imag} */,
  {32'h4236942c, 32'hc2c27fb2} /* (15, 14, 25) {real, imag} */,
  {32'hc15abdb0, 32'hc31f4ca8} /* (15, 14, 24) {real, imag} */,
  {32'hc237dc8e, 32'hc0b8ce1c} /* (15, 14, 23) {real, imag} */,
  {32'hc2a54941, 32'h42c35fd3} /* (15, 14, 22) {real, imag} */,
  {32'h42236602, 32'h4199661e} /* (15, 14, 21) {real, imag} */,
  {32'h42222ae0, 32'hc0f29704} /* (15, 14, 20) {real, imag} */,
  {32'h428505c9, 32'h425927b2} /* (15, 14, 19) {real, imag} */,
  {32'hc23751b7, 32'hc1eaf0a8} /* (15, 14, 18) {real, imag} */,
  {32'h424b9a7e, 32'h429a049d} /* (15, 14, 17) {real, imag} */,
  {32'h42043880, 32'h00000000} /* (15, 14, 16) {real, imag} */,
  {32'h424b9a7e, 32'hc29a049d} /* (15, 14, 15) {real, imag} */,
  {32'hc23751b7, 32'h41eaf0a8} /* (15, 14, 14) {real, imag} */,
  {32'h428505c9, 32'hc25927b2} /* (15, 14, 13) {real, imag} */,
  {32'h42222ae0, 32'h40f29704} /* (15, 14, 12) {real, imag} */,
  {32'h42236602, 32'hc199661e} /* (15, 14, 11) {real, imag} */,
  {32'hc2a54941, 32'hc2c35fd3} /* (15, 14, 10) {real, imag} */,
  {32'hc237dc8e, 32'h40b8ce1c} /* (15, 14, 9) {real, imag} */,
  {32'hc15abdb0, 32'h431f4ca8} /* (15, 14, 8) {real, imag} */,
  {32'h4236942c, 32'h42c27fb2} /* (15, 14, 7) {real, imag} */,
  {32'h41b8cdc8, 32'h42188bc8} /* (15, 14, 6) {real, imag} */,
  {32'h4035dc90, 32'h43128fed} /* (15, 14, 5) {real, imag} */,
  {32'hc217590c, 32'hc321be90} /* (15, 14, 4) {real, imag} */,
  {32'h43274f4e, 32'h418a35fa} /* (15, 14, 3) {real, imag} */,
  {32'h44023bfd, 32'hc2b83523} /* (15, 14, 2) {real, imag} */,
  {32'hc4a31fed, 32'hc3e1bec1} /* (15, 14, 1) {real, imag} */,
  {32'hc4289f06, 32'h00000000} /* (15, 14, 0) {real, imag} */,
  {32'hc4766b5b, 32'h43c22016} /* (15, 13, 31) {real, imag} */,
  {32'h43e35c20, 32'hc296d9af} /* (15, 13, 30) {real, imag} */,
  {32'h423aab92, 32'hc09b3f8c} /* (15, 13, 29) {real, imag} */,
  {32'hc297fdfb, 32'h4345e610} /* (15, 13, 28) {real, imag} */,
  {32'h423c4446, 32'hc172edfc} /* (15, 13, 27) {real, imag} */,
  {32'hc27c66eb, 32'hc2873398} /* (15, 13, 26) {real, imag} */,
  {32'h42b574e8, 32'hc2361449} /* (15, 13, 25) {real, imag} */,
  {32'hc07f8958, 32'hc15e0dc0} /* (15, 13, 24) {real, imag} */,
  {32'hc215359f, 32'h429d4ffa} /* (15, 13, 23) {real, imag} */,
  {32'hc2cc31b2, 32'hc28cedad} /* (15, 13, 22) {real, imag} */,
  {32'hc25aaa24, 32'hc269541c} /* (15, 13, 21) {real, imag} */,
  {32'h403f67d0, 32'h410444ec} /* (15, 13, 20) {real, imag} */,
  {32'hc20451ac, 32'h40dcd2d0} /* (15, 13, 19) {real, imag} */,
  {32'h40cb809a, 32'h420c73e3} /* (15, 13, 18) {real, imag} */,
  {32'hc2ab9034, 32'h419c6b72} /* (15, 13, 17) {real, imag} */,
  {32'hc1b8cfee, 32'h00000000} /* (15, 13, 16) {real, imag} */,
  {32'hc2ab9034, 32'hc19c6b72} /* (15, 13, 15) {real, imag} */,
  {32'h40cb809a, 32'hc20c73e3} /* (15, 13, 14) {real, imag} */,
  {32'hc20451ac, 32'hc0dcd2d0} /* (15, 13, 13) {real, imag} */,
  {32'h403f67d0, 32'hc10444ec} /* (15, 13, 12) {real, imag} */,
  {32'hc25aaa24, 32'h4269541c} /* (15, 13, 11) {real, imag} */,
  {32'hc2cc31b2, 32'h428cedad} /* (15, 13, 10) {real, imag} */,
  {32'hc215359f, 32'hc29d4ffa} /* (15, 13, 9) {real, imag} */,
  {32'hc07f8958, 32'h415e0dc0} /* (15, 13, 8) {real, imag} */,
  {32'h42b574e8, 32'h42361449} /* (15, 13, 7) {real, imag} */,
  {32'hc27c66eb, 32'h42873398} /* (15, 13, 6) {real, imag} */,
  {32'h423c4446, 32'h4172edfc} /* (15, 13, 5) {real, imag} */,
  {32'hc297fdfb, 32'hc345e610} /* (15, 13, 4) {real, imag} */,
  {32'h423aab92, 32'h409b3f8c} /* (15, 13, 3) {real, imag} */,
  {32'h43e35c20, 32'h4296d9af} /* (15, 13, 2) {real, imag} */,
  {32'hc4766b5b, 32'hc3c22016} /* (15, 13, 1) {real, imag} */,
  {32'hc3f487ac, 32'h00000000} /* (15, 13, 0) {real, imag} */,
  {32'hc451fcc1, 32'h437ebcdc} /* (15, 12, 31) {real, imag} */,
  {32'h43b28bbe, 32'h403c3690} /* (15, 12, 30) {real, imag} */,
  {32'h42529a5a, 32'h4147cb48} /* (15, 12, 29) {real, imag} */,
  {32'hc341a85a, 32'h4310c1cc} /* (15, 12, 28) {real, imag} */,
  {32'h429f17e1, 32'hc2dbc7eb} /* (15, 12, 27) {real, imag} */,
  {32'h4303a618, 32'h432bc639} /* (15, 12, 26) {real, imag} */,
  {32'hc2be1398, 32'hc0b276c0} /* (15, 12, 25) {real, imag} */,
  {32'h42d17254, 32'h4147911c} /* (15, 12, 24) {real, imag} */,
  {32'hc2a771b0, 32'hc2158670} /* (15, 12, 23) {real, imag} */,
  {32'h4215e302, 32'hc01df4ee} /* (15, 12, 22) {real, imag} */,
  {32'h4134c3f7, 32'hc1e4db50} /* (15, 12, 21) {real, imag} */,
  {32'hc29a8674, 32'h40a6bc02} /* (15, 12, 20) {real, imag} */,
  {32'hc2a79299, 32'hc2802386} /* (15, 12, 19) {real, imag} */,
  {32'h4292be4e, 32'h420f1136} /* (15, 12, 18) {real, imag} */,
  {32'h4174c267, 32'h420bb792} /* (15, 12, 17) {real, imag} */,
  {32'h403db4a8, 32'h00000000} /* (15, 12, 16) {real, imag} */,
  {32'h4174c267, 32'hc20bb792} /* (15, 12, 15) {real, imag} */,
  {32'h4292be4e, 32'hc20f1136} /* (15, 12, 14) {real, imag} */,
  {32'hc2a79299, 32'h42802386} /* (15, 12, 13) {real, imag} */,
  {32'hc29a8674, 32'hc0a6bc02} /* (15, 12, 12) {real, imag} */,
  {32'h4134c3f7, 32'h41e4db50} /* (15, 12, 11) {real, imag} */,
  {32'h4215e302, 32'h401df4ee} /* (15, 12, 10) {real, imag} */,
  {32'hc2a771b0, 32'h42158670} /* (15, 12, 9) {real, imag} */,
  {32'h42d17254, 32'hc147911c} /* (15, 12, 8) {real, imag} */,
  {32'hc2be1398, 32'h40b276c0} /* (15, 12, 7) {real, imag} */,
  {32'h4303a618, 32'hc32bc639} /* (15, 12, 6) {real, imag} */,
  {32'h429f17e1, 32'h42dbc7eb} /* (15, 12, 5) {real, imag} */,
  {32'hc341a85a, 32'hc310c1cc} /* (15, 12, 4) {real, imag} */,
  {32'h42529a5a, 32'hc147cb48} /* (15, 12, 3) {real, imag} */,
  {32'h43b28bbe, 32'hc03c3690} /* (15, 12, 2) {real, imag} */,
  {32'hc451fcc1, 32'hc37ebcdc} /* (15, 12, 1) {real, imag} */,
  {32'h4167c160, 32'h00000000} /* (15, 12, 0) {real, imag} */,
  {32'hc40f5e10, 32'h431d23a7} /* (15, 11, 31) {real, imag} */,
  {32'h43b9b12e, 32'h42ace6e6} /* (15, 11, 30) {real, imag} */,
  {32'h4203712c, 32'hc1bae330} /* (15, 11, 29) {real, imag} */,
  {32'hc30dad72, 32'h42d87d82} /* (15, 11, 28) {real, imag} */,
  {32'h42dadd33, 32'hc2a2bc13} /* (15, 11, 27) {real, imag} */,
  {32'h428b1397, 32'hc294ce8c} /* (15, 11, 26) {real, imag} */,
  {32'hc319677d, 32'h416a1158} /* (15, 11, 25) {real, imag} */,
  {32'hc187d3b8, 32'hc216c68c} /* (15, 11, 24) {real, imag} */,
  {32'h426b72cb, 32'hc2b1ffd6} /* (15, 11, 23) {real, imag} */,
  {32'hc2c8cd01, 32'hc23c3087} /* (15, 11, 22) {real, imag} */,
  {32'hc1a11f72, 32'h421e4c4c} /* (15, 11, 21) {real, imag} */,
  {32'h42b8bd20, 32'h4296e12d} /* (15, 11, 20) {real, imag} */,
  {32'hc2a320db, 32'hc264de8b} /* (15, 11, 19) {real, imag} */,
  {32'hc1c26082, 32'hc2862c5c} /* (15, 11, 18) {real, imag} */,
  {32'h41464444, 32'h42d11a84} /* (15, 11, 17) {real, imag} */,
  {32'h41dabfa0, 32'h00000000} /* (15, 11, 16) {real, imag} */,
  {32'h41464444, 32'hc2d11a84} /* (15, 11, 15) {real, imag} */,
  {32'hc1c26082, 32'h42862c5c} /* (15, 11, 14) {real, imag} */,
  {32'hc2a320db, 32'h4264de8b} /* (15, 11, 13) {real, imag} */,
  {32'h42b8bd20, 32'hc296e12d} /* (15, 11, 12) {real, imag} */,
  {32'hc1a11f72, 32'hc21e4c4c} /* (15, 11, 11) {real, imag} */,
  {32'hc2c8cd01, 32'h423c3087} /* (15, 11, 10) {real, imag} */,
  {32'h426b72cb, 32'h42b1ffd6} /* (15, 11, 9) {real, imag} */,
  {32'hc187d3b8, 32'h4216c68c} /* (15, 11, 8) {real, imag} */,
  {32'hc319677d, 32'hc16a1158} /* (15, 11, 7) {real, imag} */,
  {32'h428b1397, 32'h4294ce8c} /* (15, 11, 6) {real, imag} */,
  {32'h42dadd33, 32'h42a2bc13} /* (15, 11, 5) {real, imag} */,
  {32'hc30dad72, 32'hc2d87d82} /* (15, 11, 4) {real, imag} */,
  {32'h4203712c, 32'h41bae330} /* (15, 11, 3) {real, imag} */,
  {32'h43b9b12e, 32'hc2ace6e6} /* (15, 11, 2) {real, imag} */,
  {32'hc40f5e10, 32'hc31d23a7} /* (15, 11, 1) {real, imag} */,
  {32'h43caf990, 32'h00000000} /* (15, 11, 0) {real, imag} */,
  {32'h43163062, 32'h42c5dec9} /* (15, 10, 31) {real, imag} */,
  {32'h42e017a2, 32'h430bf050} /* (15, 10, 30) {real, imag} */,
  {32'hc21be906, 32'hc2a76b74} /* (15, 10, 29) {real, imag} */,
  {32'hc2787f8f, 32'hc1c015b8} /* (15, 10, 28) {real, imag} */,
  {32'hc24dbeaa, 32'h42902aa8} /* (15, 10, 27) {real, imag} */,
  {32'h41b13544, 32'h4212ad5d} /* (15, 10, 26) {real, imag} */,
  {32'hc2810f4e, 32'hc2a89853} /* (15, 10, 25) {real, imag} */,
  {32'hc30d4e1f, 32'h432e2746} /* (15, 10, 24) {real, imag} */,
  {32'h4281574c, 32'h41b596dc} /* (15, 10, 23) {real, imag} */,
  {32'hc261fa1c, 32'hc213b9dc} /* (15, 10, 22) {real, imag} */,
  {32'hc15e7ea9, 32'hc29594ac} /* (15, 10, 21) {real, imag} */,
  {32'h428d9ed0, 32'h41e4b978} /* (15, 10, 20) {real, imag} */,
  {32'h43053681, 32'hc2437082} /* (15, 10, 19) {real, imag} */,
  {32'h41e7ff9b, 32'hc182a06e} /* (15, 10, 18) {real, imag} */,
  {32'hc2496850, 32'h4310693f} /* (15, 10, 17) {real, imag} */,
  {32'h42973f44, 32'h00000000} /* (15, 10, 16) {real, imag} */,
  {32'hc2496850, 32'hc310693f} /* (15, 10, 15) {real, imag} */,
  {32'h41e7ff9b, 32'h4182a06e} /* (15, 10, 14) {real, imag} */,
  {32'h43053681, 32'h42437082} /* (15, 10, 13) {real, imag} */,
  {32'h428d9ed0, 32'hc1e4b978} /* (15, 10, 12) {real, imag} */,
  {32'hc15e7ea9, 32'h429594ac} /* (15, 10, 11) {real, imag} */,
  {32'hc261fa1c, 32'h4213b9dc} /* (15, 10, 10) {real, imag} */,
  {32'h4281574c, 32'hc1b596dc} /* (15, 10, 9) {real, imag} */,
  {32'hc30d4e1f, 32'hc32e2746} /* (15, 10, 8) {real, imag} */,
  {32'hc2810f4e, 32'h42a89853} /* (15, 10, 7) {real, imag} */,
  {32'h41b13544, 32'hc212ad5d} /* (15, 10, 6) {real, imag} */,
  {32'hc24dbeaa, 32'hc2902aa8} /* (15, 10, 5) {real, imag} */,
  {32'hc2787f8f, 32'h41c015b8} /* (15, 10, 4) {real, imag} */,
  {32'hc21be906, 32'h42a76b74} /* (15, 10, 3) {real, imag} */,
  {32'h42e017a2, 32'hc30bf050} /* (15, 10, 2) {real, imag} */,
  {32'h43163062, 32'hc2c5dec9} /* (15, 10, 1) {real, imag} */,
  {32'h4445c425, 32'h00000000} /* (15, 10, 0) {real, imag} */,
  {32'h43d0f1d8, 32'hc23af246} /* (15, 9, 31) {real, imag} */,
  {32'hc2d17a6a, 32'h433ae886} /* (15, 9, 30) {real, imag} */,
  {32'hc2f7c778, 32'h425282a0} /* (15, 9, 29) {real, imag} */,
  {32'hc26ec624, 32'hc1ae48fc} /* (15, 9, 28) {real, imag} */,
  {32'hc2fa9e31, 32'hc16c9bc6} /* (15, 9, 27) {real, imag} */,
  {32'h4291fc58, 32'h4311d05a} /* (15, 9, 26) {real, imag} */,
  {32'h424304fc, 32'hc299b97d} /* (15, 9, 25) {real, imag} */,
  {32'hc04892e8, 32'h426ead09} /* (15, 9, 24) {real, imag} */,
  {32'hc27ad7df, 32'hc0d2d0ad} /* (15, 9, 23) {real, imag} */,
  {32'h42dff422, 32'hc29a8e7a} /* (15, 9, 22) {real, imag} */,
  {32'hc1d24988, 32'hc2710b9a} /* (15, 9, 21) {real, imag} */,
  {32'hc00f6cb8, 32'h42a16a9f} /* (15, 9, 20) {real, imag} */,
  {32'hc2fdc688, 32'hc1849f40} /* (15, 9, 19) {real, imag} */,
  {32'h41e07239, 32'h420c52b7} /* (15, 9, 18) {real, imag} */,
  {32'hc2922756, 32'h41e11d5c} /* (15, 9, 17) {real, imag} */,
  {32'h42d920fe, 32'h00000000} /* (15, 9, 16) {real, imag} */,
  {32'hc2922756, 32'hc1e11d5c} /* (15, 9, 15) {real, imag} */,
  {32'h41e07239, 32'hc20c52b7} /* (15, 9, 14) {real, imag} */,
  {32'hc2fdc688, 32'h41849f40} /* (15, 9, 13) {real, imag} */,
  {32'hc00f6cb8, 32'hc2a16a9f} /* (15, 9, 12) {real, imag} */,
  {32'hc1d24988, 32'h42710b9a} /* (15, 9, 11) {real, imag} */,
  {32'h42dff422, 32'h429a8e7a} /* (15, 9, 10) {real, imag} */,
  {32'hc27ad7df, 32'h40d2d0ad} /* (15, 9, 9) {real, imag} */,
  {32'hc04892e8, 32'hc26ead09} /* (15, 9, 8) {real, imag} */,
  {32'h424304fc, 32'h4299b97d} /* (15, 9, 7) {real, imag} */,
  {32'h4291fc58, 32'hc311d05a} /* (15, 9, 6) {real, imag} */,
  {32'hc2fa9e31, 32'h416c9bc6} /* (15, 9, 5) {real, imag} */,
  {32'hc26ec624, 32'h41ae48fc} /* (15, 9, 4) {real, imag} */,
  {32'hc2f7c778, 32'hc25282a0} /* (15, 9, 3) {real, imag} */,
  {32'hc2d17a6a, 32'hc33ae886} /* (15, 9, 2) {real, imag} */,
  {32'h43d0f1d8, 32'h423af246} /* (15, 9, 1) {real, imag} */,
  {32'h447aac80, 32'h00000000} /* (15, 9, 0) {real, imag} */,
  {32'h43ea8a56, 32'hc32f7f8f} /* (15, 8, 31) {real, imag} */,
  {32'hc3937051, 32'h4365a604} /* (15, 8, 30) {real, imag} */,
  {32'hc327e8ee, 32'hc1a5f018} /* (15, 8, 29) {real, imag} */,
  {32'hc17c60ba, 32'hc2d9b348} /* (15, 8, 28) {real, imag} */,
  {32'hc2e45732, 32'h42b4d965} /* (15, 8, 27) {real, imag} */,
  {32'h42c06e56, 32'hc1bba3ba} /* (15, 8, 26) {real, imag} */,
  {32'hc1fe6ff9, 32'hc1d90afc} /* (15, 8, 25) {real, imag} */,
  {32'hc2c510a1, 32'h42cf688e} /* (15, 8, 24) {real, imag} */,
  {32'hc22189cd, 32'hc299e2e8} /* (15, 8, 23) {real, imag} */,
  {32'h42a1ba26, 32'h4221442a} /* (15, 8, 22) {real, imag} */,
  {32'h4291ed3a, 32'h42eb50af} /* (15, 8, 21) {real, imag} */,
  {32'h4302d50e, 32'h42acda66} /* (15, 8, 20) {real, imag} */,
  {32'hc2ae1991, 32'hc00ca80c} /* (15, 8, 19) {real, imag} */,
  {32'hc187b383, 32'h418b87b9} /* (15, 8, 18) {real, imag} */,
  {32'h42b922fa, 32'hc2ae0075} /* (15, 8, 17) {real, imag} */,
  {32'h426eec10, 32'h00000000} /* (15, 8, 16) {real, imag} */,
  {32'h42b922fa, 32'h42ae0075} /* (15, 8, 15) {real, imag} */,
  {32'hc187b383, 32'hc18b87b9} /* (15, 8, 14) {real, imag} */,
  {32'hc2ae1991, 32'h400ca80c} /* (15, 8, 13) {real, imag} */,
  {32'h4302d50e, 32'hc2acda66} /* (15, 8, 12) {real, imag} */,
  {32'h4291ed3a, 32'hc2eb50af} /* (15, 8, 11) {real, imag} */,
  {32'h42a1ba26, 32'hc221442a} /* (15, 8, 10) {real, imag} */,
  {32'hc22189cd, 32'h4299e2e8} /* (15, 8, 9) {real, imag} */,
  {32'hc2c510a1, 32'hc2cf688e} /* (15, 8, 8) {real, imag} */,
  {32'hc1fe6ff9, 32'h41d90afc} /* (15, 8, 7) {real, imag} */,
  {32'h42c06e56, 32'h41bba3ba} /* (15, 8, 6) {real, imag} */,
  {32'hc2e45732, 32'hc2b4d965} /* (15, 8, 5) {real, imag} */,
  {32'hc17c60ba, 32'h42d9b348} /* (15, 8, 4) {real, imag} */,
  {32'hc327e8ee, 32'h41a5f018} /* (15, 8, 3) {real, imag} */,
  {32'hc3937051, 32'hc365a604} /* (15, 8, 2) {real, imag} */,
  {32'h43ea8a56, 32'h432f7f8f} /* (15, 8, 1) {real, imag} */,
  {32'h4481d877, 32'h00000000} /* (15, 8, 0) {real, imag} */,
  {32'h44137dd2, 32'hc3035fe4} /* (15, 7, 31) {real, imag} */,
  {32'hc3a0f27e, 32'h433455dc} /* (15, 7, 30) {real, imag} */,
  {32'hc27e14a8, 32'hc26efbda} /* (15, 7, 29) {real, imag} */,
  {32'h4261afb4, 32'hc3034f0c} /* (15, 7, 28) {real, imag} */,
  {32'hc31ca6c5, 32'hc1a0dc54} /* (15, 7, 27) {real, imag} */,
  {32'h4263490f, 32'h3f4ef7e0} /* (15, 7, 26) {real, imag} */,
  {32'hc0eb5e30, 32'hc2362e38} /* (15, 7, 25) {real, imag} */,
  {32'hc23ea9ec, 32'h42576d4f} /* (15, 7, 24) {real, imag} */,
  {32'h42bae2b6, 32'h42180c82} /* (15, 7, 23) {real, imag} */,
  {32'hc18170b7, 32'h4296fe9e} /* (15, 7, 22) {real, imag} */,
  {32'hc2284fa0, 32'hc24536c0} /* (15, 7, 21) {real, imag} */,
  {32'h41e66beb, 32'hc17d5d1c} /* (15, 7, 20) {real, imag} */,
  {32'h427663de, 32'h41e4d6f0} /* (15, 7, 19) {real, imag} */,
  {32'hc28762ef, 32'h42495775} /* (15, 7, 18) {real, imag} */,
  {32'hc1aab788, 32'hc1aa1479} /* (15, 7, 17) {real, imag} */,
  {32'hc2606c24, 32'h00000000} /* (15, 7, 16) {real, imag} */,
  {32'hc1aab788, 32'h41aa1479} /* (15, 7, 15) {real, imag} */,
  {32'hc28762ef, 32'hc2495775} /* (15, 7, 14) {real, imag} */,
  {32'h427663de, 32'hc1e4d6f0} /* (15, 7, 13) {real, imag} */,
  {32'h41e66beb, 32'h417d5d1c} /* (15, 7, 12) {real, imag} */,
  {32'hc2284fa0, 32'h424536c0} /* (15, 7, 11) {real, imag} */,
  {32'hc18170b7, 32'hc296fe9e} /* (15, 7, 10) {real, imag} */,
  {32'h42bae2b6, 32'hc2180c82} /* (15, 7, 9) {real, imag} */,
  {32'hc23ea9ec, 32'hc2576d4f} /* (15, 7, 8) {real, imag} */,
  {32'hc0eb5e30, 32'h42362e38} /* (15, 7, 7) {real, imag} */,
  {32'h4263490f, 32'hbf4ef7e0} /* (15, 7, 6) {real, imag} */,
  {32'hc31ca6c5, 32'h41a0dc54} /* (15, 7, 5) {real, imag} */,
  {32'h4261afb4, 32'h43034f0c} /* (15, 7, 4) {real, imag} */,
  {32'hc27e14a8, 32'h426efbda} /* (15, 7, 3) {real, imag} */,
  {32'hc3a0f27e, 32'hc33455dc} /* (15, 7, 2) {real, imag} */,
  {32'h44137dd2, 32'h43035fe4} /* (15, 7, 1) {real, imag} */,
  {32'h448fe642, 32'h00000000} /* (15, 7, 0) {real, imag} */,
  {32'h44060ce9, 32'hc37057ec} /* (15, 6, 31) {real, imag} */,
  {32'hc3b1347e, 32'h435852ba} /* (15, 6, 30) {real, imag} */,
  {32'hbfc980b0, 32'h42ffa988} /* (15, 6, 29) {real, imag} */,
  {32'h41b4af7a, 32'hc2b5d246} /* (15, 6, 28) {real, imag} */,
  {32'hc289fbfb, 32'h417dba70} /* (15, 6, 27) {real, imag} */,
  {32'h42774781, 32'hc28ae9f4} /* (15, 6, 26) {real, imag} */,
  {32'h41e45b5c, 32'hc206ea9a} /* (15, 6, 25) {real, imag} */,
  {32'hc216b851, 32'h41957ade} /* (15, 6, 24) {real, imag} */,
  {32'hc14695c8, 32'h4225ae11} /* (15, 6, 23) {real, imag} */,
  {32'hc250111c, 32'h41a19f42} /* (15, 6, 22) {real, imag} */,
  {32'hc1e9ad49, 32'h41434d28} /* (15, 6, 21) {real, imag} */,
  {32'h4213c718, 32'hc2825eaa} /* (15, 6, 20) {real, imag} */,
  {32'hc225cc6e, 32'h42300829} /* (15, 6, 19) {real, imag} */,
  {32'hc208073c, 32'h427645b1} /* (15, 6, 18) {real, imag} */,
  {32'h423acaec, 32'h413fb2b4} /* (15, 6, 17) {real, imag} */,
  {32'h4227adfd, 32'h00000000} /* (15, 6, 16) {real, imag} */,
  {32'h423acaec, 32'hc13fb2b4} /* (15, 6, 15) {real, imag} */,
  {32'hc208073c, 32'hc27645b1} /* (15, 6, 14) {real, imag} */,
  {32'hc225cc6e, 32'hc2300829} /* (15, 6, 13) {real, imag} */,
  {32'h4213c718, 32'h42825eaa} /* (15, 6, 12) {real, imag} */,
  {32'hc1e9ad49, 32'hc1434d28} /* (15, 6, 11) {real, imag} */,
  {32'hc250111c, 32'hc1a19f42} /* (15, 6, 10) {real, imag} */,
  {32'hc14695c8, 32'hc225ae11} /* (15, 6, 9) {real, imag} */,
  {32'hc216b851, 32'hc1957ade} /* (15, 6, 8) {real, imag} */,
  {32'h41e45b5c, 32'h4206ea9a} /* (15, 6, 7) {real, imag} */,
  {32'h42774781, 32'h428ae9f4} /* (15, 6, 6) {real, imag} */,
  {32'hc289fbfb, 32'hc17dba70} /* (15, 6, 5) {real, imag} */,
  {32'h41b4af7a, 32'h42b5d246} /* (15, 6, 4) {real, imag} */,
  {32'hbfc980b0, 32'hc2ffa988} /* (15, 6, 3) {real, imag} */,
  {32'hc3b1347e, 32'hc35852ba} /* (15, 6, 2) {real, imag} */,
  {32'h44060ce9, 32'h437057ec} /* (15, 6, 1) {real, imag} */,
  {32'h448a4351, 32'h00000000} /* (15, 6, 0) {real, imag} */,
  {32'h4424e6d7, 32'hc4141149} /* (15, 5, 31) {real, imag} */,
  {32'hc337133d, 32'h4384f25b} /* (15, 5, 30) {real, imag} */,
  {32'hc325f50c, 32'h42ebef97} /* (15, 5, 29) {real, imag} */,
  {32'hc2a4c2fd, 32'hc2d99c5d} /* (15, 5, 28) {real, imag} */,
  {32'hc2a447d6, 32'hbfec4080} /* (15, 5, 27) {real, imag} */,
  {32'hc2096878, 32'hc2a30369} /* (15, 5, 26) {real, imag} */,
  {32'h42dc91c2, 32'hc1252fe0} /* (15, 5, 25) {real, imag} */,
  {32'h42d32b94, 32'h423b2ec8} /* (15, 5, 24) {real, imag} */,
  {32'hc2efb6cc, 32'hc1b6148c} /* (15, 5, 23) {real, imag} */,
  {32'hc246c526, 32'h41c288a6} /* (15, 5, 22) {real, imag} */,
  {32'hc1e7b32e, 32'h42abbae6} /* (15, 5, 21) {real, imag} */,
  {32'hc1b3c7f6, 32'h426ad658} /* (15, 5, 20) {real, imag} */,
  {32'hc2e5034a, 32'h4284d6fb} /* (15, 5, 19) {real, imag} */,
  {32'hc0d5fa80, 32'hc2e99f8f} /* (15, 5, 18) {real, imag} */,
  {32'h42a44032, 32'h42826ab7} /* (15, 5, 17) {real, imag} */,
  {32'h42e5db73, 32'h00000000} /* (15, 5, 16) {real, imag} */,
  {32'h42a44032, 32'hc2826ab7} /* (15, 5, 15) {real, imag} */,
  {32'hc0d5fa80, 32'h42e99f8f} /* (15, 5, 14) {real, imag} */,
  {32'hc2e5034a, 32'hc284d6fb} /* (15, 5, 13) {real, imag} */,
  {32'hc1b3c7f6, 32'hc26ad658} /* (15, 5, 12) {real, imag} */,
  {32'hc1e7b32e, 32'hc2abbae6} /* (15, 5, 11) {real, imag} */,
  {32'hc246c526, 32'hc1c288a6} /* (15, 5, 10) {real, imag} */,
  {32'hc2efb6cc, 32'h41b6148c} /* (15, 5, 9) {real, imag} */,
  {32'h42d32b94, 32'hc23b2ec8} /* (15, 5, 8) {real, imag} */,
  {32'h42dc91c2, 32'h41252fe0} /* (15, 5, 7) {real, imag} */,
  {32'hc2096878, 32'h42a30369} /* (15, 5, 6) {real, imag} */,
  {32'hc2a447d6, 32'h3fec4080} /* (15, 5, 5) {real, imag} */,
  {32'hc2a4c2fd, 32'h42d99c5d} /* (15, 5, 4) {real, imag} */,
  {32'hc325f50c, 32'hc2ebef97} /* (15, 5, 3) {real, imag} */,
  {32'hc337133d, 32'hc384f25b} /* (15, 5, 2) {real, imag} */,
  {32'h4424e6d7, 32'h44141149} /* (15, 5, 1) {real, imag} */,
  {32'h4485f083, 32'h00000000} /* (15, 5, 0) {real, imag} */,
  {32'h4410ca53, 32'hc44eab07} /* (15, 4, 31) {real, imag} */,
  {32'hc20ee558, 32'h43921ca6} /* (15, 4, 30) {real, imag} */,
  {32'hc2547fc9, 32'h4308b5e3} /* (15, 4, 29) {real, imag} */,
  {32'hc2d688c0, 32'h42079968} /* (15, 4, 28) {real, imag} */,
  {32'hc3005005, 32'hc1350222} /* (15, 4, 27) {real, imag} */,
  {32'h40dc2770, 32'hc0c7a684} /* (15, 4, 26) {real, imag} */,
  {32'h41d00a84, 32'hc19a8278} /* (15, 4, 25) {real, imag} */,
  {32'h422739f1, 32'h426931eb} /* (15, 4, 24) {real, imag} */,
  {32'hc16e6130, 32'hc2c39890} /* (15, 4, 23) {real, imag} */,
  {32'h41f685be, 32'h41850cd8} /* (15, 4, 22) {real, imag} */,
  {32'h41ee019c, 32'h42b64972} /* (15, 4, 21) {real, imag} */,
  {32'hc18d19ba, 32'h41908a67} /* (15, 4, 20) {real, imag} */,
  {32'h426944de, 32'hc28854b8} /* (15, 4, 19) {real, imag} */,
  {32'h40176938, 32'h42999764} /* (15, 4, 18) {real, imag} */,
  {32'hc27b7d3b, 32'hc008f426} /* (15, 4, 17) {real, imag} */,
  {32'h42c8a3b2, 32'h00000000} /* (15, 4, 16) {real, imag} */,
  {32'hc27b7d3b, 32'h4008f426} /* (15, 4, 15) {real, imag} */,
  {32'h40176938, 32'hc2999764} /* (15, 4, 14) {real, imag} */,
  {32'h426944de, 32'h428854b8} /* (15, 4, 13) {real, imag} */,
  {32'hc18d19ba, 32'hc1908a67} /* (15, 4, 12) {real, imag} */,
  {32'h41ee019c, 32'hc2b64972} /* (15, 4, 11) {real, imag} */,
  {32'h41f685be, 32'hc1850cd8} /* (15, 4, 10) {real, imag} */,
  {32'hc16e6130, 32'h42c39890} /* (15, 4, 9) {real, imag} */,
  {32'h422739f1, 32'hc26931eb} /* (15, 4, 8) {real, imag} */,
  {32'h41d00a84, 32'h419a8278} /* (15, 4, 7) {real, imag} */,
  {32'h40dc2770, 32'h40c7a684} /* (15, 4, 6) {real, imag} */,
  {32'hc3005005, 32'h41350222} /* (15, 4, 5) {real, imag} */,
  {32'hc2d688c0, 32'hc2079968} /* (15, 4, 4) {real, imag} */,
  {32'hc2547fc9, 32'hc308b5e3} /* (15, 4, 3) {real, imag} */,
  {32'hc20ee558, 32'hc3921ca6} /* (15, 4, 2) {real, imag} */,
  {32'h4410ca53, 32'h444eab07} /* (15, 4, 1) {real, imag} */,
  {32'h4494a8bc, 32'h00000000} /* (15, 4, 0) {real, imag} */,
  {32'h4428cb0d, 32'hc43f1f3a} /* (15, 3, 31) {real, imag} */,
  {32'hc25af77c, 32'h43bc6983} /* (15, 3, 30) {real, imag} */,
  {32'hc262d89c, 32'h42927d4c} /* (15, 3, 29) {real, imag} */,
  {32'hc32bb559, 32'h4281c4ae} /* (15, 3, 28) {real, imag} */,
  {32'hc2e39dda, 32'hc30390f3} /* (15, 3, 27) {real, imag} */,
  {32'h425bd4dd, 32'hc1f9232b} /* (15, 3, 26) {real, imag} */,
  {32'h421a738d, 32'hc3030a95} /* (15, 3, 25) {real, imag} */,
  {32'h42083604, 32'hc0efa084} /* (15, 3, 24) {real, imag} */,
  {32'h4258fa06, 32'h419b7aae} /* (15, 3, 23) {real, imag} */,
  {32'h4288ba3f, 32'h4245a270} /* (15, 3, 22) {real, imag} */,
  {32'hc1f50ca4, 32'hc114222e} /* (15, 3, 21) {real, imag} */,
  {32'h42678990, 32'hc1875a32} /* (15, 3, 20) {real, imag} */,
  {32'hc22777b0, 32'h42256761} /* (15, 3, 19) {real, imag} */,
  {32'hc170ebc0, 32'h41b3fda2} /* (15, 3, 18) {real, imag} */,
  {32'hc2901ea2, 32'h42946184} /* (15, 3, 17) {real, imag} */,
  {32'h42a2185c, 32'h00000000} /* (15, 3, 16) {real, imag} */,
  {32'hc2901ea2, 32'hc2946184} /* (15, 3, 15) {real, imag} */,
  {32'hc170ebc0, 32'hc1b3fda2} /* (15, 3, 14) {real, imag} */,
  {32'hc22777b0, 32'hc2256761} /* (15, 3, 13) {real, imag} */,
  {32'h42678990, 32'h41875a32} /* (15, 3, 12) {real, imag} */,
  {32'hc1f50ca4, 32'h4114222e} /* (15, 3, 11) {real, imag} */,
  {32'h4288ba3f, 32'hc245a270} /* (15, 3, 10) {real, imag} */,
  {32'h4258fa06, 32'hc19b7aae} /* (15, 3, 9) {real, imag} */,
  {32'h42083604, 32'h40efa084} /* (15, 3, 8) {real, imag} */,
  {32'h421a738d, 32'h43030a95} /* (15, 3, 7) {real, imag} */,
  {32'h425bd4dd, 32'h41f9232b} /* (15, 3, 6) {real, imag} */,
  {32'hc2e39dda, 32'h430390f3} /* (15, 3, 5) {real, imag} */,
  {32'hc32bb559, 32'hc281c4ae} /* (15, 3, 4) {real, imag} */,
  {32'hc262d89c, 32'hc2927d4c} /* (15, 3, 3) {real, imag} */,
  {32'hc25af77c, 32'hc3bc6983} /* (15, 3, 2) {real, imag} */,
  {32'h4428cb0d, 32'h443f1f3a} /* (15, 3, 1) {real, imag} */,
  {32'h44a3c3dd, 32'h00000000} /* (15, 3, 0) {real, imag} */,
  {32'h4422520b, 32'hc4421e5b} /* (15, 2, 31) {real, imag} */,
  {32'h429756b6, 32'h439c73a6} /* (15, 2, 30) {real, imag} */,
  {32'hc317081e, 32'h41085654} /* (15, 2, 29) {real, imag} */,
  {32'hc1d6b132, 32'h42473dfc} /* (15, 2, 28) {real, imag} */,
  {32'hc322c92e, 32'hc2bf9454} /* (15, 2, 27) {real, imag} */,
  {32'hc0a0b520, 32'hbfadc9f0} /* (15, 2, 26) {real, imag} */,
  {32'hc1b596c4, 32'hc222d230} /* (15, 2, 25) {real, imag} */,
  {32'h42784639, 32'h41164fe6} /* (15, 2, 24) {real, imag} */,
  {32'hc2fffa53, 32'h417ef31c} /* (15, 2, 23) {real, imag} */,
  {32'h3fef9380, 32'h419fd42c} /* (15, 2, 22) {real, imag} */,
  {32'hc2a0503d, 32'h409a5884} /* (15, 2, 21) {real, imag} */,
  {32'h42733742, 32'hc1d29489} /* (15, 2, 20) {real, imag} */,
  {32'h3f9f7270, 32'h4056fe00} /* (15, 2, 19) {real, imag} */,
  {32'h426326e0, 32'h42d22cc1} /* (15, 2, 18) {real, imag} */,
  {32'h420ef6c0, 32'h40ff9da0} /* (15, 2, 17) {real, imag} */,
  {32'h42b04fd6, 32'h00000000} /* (15, 2, 16) {real, imag} */,
  {32'h420ef6c0, 32'hc0ff9da0} /* (15, 2, 15) {real, imag} */,
  {32'h426326e0, 32'hc2d22cc1} /* (15, 2, 14) {real, imag} */,
  {32'h3f9f7270, 32'hc056fe00} /* (15, 2, 13) {real, imag} */,
  {32'h42733742, 32'h41d29489} /* (15, 2, 12) {real, imag} */,
  {32'hc2a0503d, 32'hc09a5884} /* (15, 2, 11) {real, imag} */,
  {32'h3fef9380, 32'hc19fd42c} /* (15, 2, 10) {real, imag} */,
  {32'hc2fffa53, 32'hc17ef31c} /* (15, 2, 9) {real, imag} */,
  {32'h42784639, 32'hc1164fe6} /* (15, 2, 8) {real, imag} */,
  {32'hc1b596c4, 32'h4222d230} /* (15, 2, 7) {real, imag} */,
  {32'hc0a0b520, 32'h3fadc9f0} /* (15, 2, 6) {real, imag} */,
  {32'hc322c92e, 32'h42bf9454} /* (15, 2, 5) {real, imag} */,
  {32'hc1d6b132, 32'hc2473dfc} /* (15, 2, 4) {real, imag} */,
  {32'hc317081e, 32'hc1085654} /* (15, 2, 3) {real, imag} */,
  {32'h429756b6, 32'hc39c73a6} /* (15, 2, 2) {real, imag} */,
  {32'h4422520b, 32'h44421e5b} /* (15, 2, 1) {real, imag} */,
  {32'h449b8f6d, 32'h00000000} /* (15, 2, 0) {real, imag} */,
  {32'h4408c6f7, 32'hc46a3331} /* (15, 1, 31) {real, imag} */,
  {32'h42a58a96, 32'h43447fc8} /* (15, 1, 30) {real, imag} */,
  {32'h4200682f, 32'h42643695} /* (15, 1, 29) {real, imag} */,
  {32'hc29068c2, 32'h42b01261} /* (15, 1, 28) {real, imag} */,
  {32'hc2d37c65, 32'h421677e2} /* (15, 1, 27) {real, imag} */,
  {32'hc236310b, 32'h42bb7822} /* (15, 1, 26) {real, imag} */,
  {32'hc29373e8, 32'hc2a725a4} /* (15, 1, 25) {real, imag} */,
  {32'h4228fe27, 32'hc1a03e8a} /* (15, 1, 24) {real, imag} */,
  {32'hc2858cb3, 32'h4089adfc} /* (15, 1, 23) {real, imag} */,
  {32'h4209faca, 32'h42801ea7} /* (15, 1, 22) {real, imag} */,
  {32'hc2d97192, 32'hc1ae0db7} /* (15, 1, 21) {real, imag} */,
  {32'hc22d726f, 32'h42834c56} /* (15, 1, 20) {real, imag} */,
  {32'h419afe26, 32'hc1c20579} /* (15, 1, 19) {real, imag} */,
  {32'h3f9048a8, 32'hc20ef7dd} /* (15, 1, 18) {real, imag} */,
  {32'h42024cdc, 32'h4117a3e1} /* (15, 1, 17) {real, imag} */,
  {32'hc2602828, 32'h00000000} /* (15, 1, 16) {real, imag} */,
  {32'h42024cdc, 32'hc117a3e1} /* (15, 1, 15) {real, imag} */,
  {32'h3f9048a8, 32'h420ef7dd} /* (15, 1, 14) {real, imag} */,
  {32'h419afe26, 32'h41c20579} /* (15, 1, 13) {real, imag} */,
  {32'hc22d726f, 32'hc2834c56} /* (15, 1, 12) {real, imag} */,
  {32'hc2d97192, 32'h41ae0db7} /* (15, 1, 11) {real, imag} */,
  {32'h4209faca, 32'hc2801ea7} /* (15, 1, 10) {real, imag} */,
  {32'hc2858cb3, 32'hc089adfc} /* (15, 1, 9) {real, imag} */,
  {32'h4228fe27, 32'h41a03e8a} /* (15, 1, 8) {real, imag} */,
  {32'hc29373e8, 32'h42a725a4} /* (15, 1, 7) {real, imag} */,
  {32'hc236310b, 32'hc2bb7822} /* (15, 1, 6) {real, imag} */,
  {32'hc2d37c65, 32'hc21677e2} /* (15, 1, 5) {real, imag} */,
  {32'hc29068c2, 32'hc2b01261} /* (15, 1, 4) {real, imag} */,
  {32'h4200682f, 32'hc2643695} /* (15, 1, 3) {real, imag} */,
  {32'h42a58a96, 32'hc3447fc8} /* (15, 1, 2) {real, imag} */,
  {32'h4408c6f7, 32'h446a3331} /* (15, 1, 1) {real, imag} */,
  {32'h444ec941, 32'h00000000} /* (15, 1, 0) {real, imag} */,
  {32'h4415afcb, 32'hc42b896b} /* (15, 0, 31) {real, imag} */,
  {32'hc1f9e1d0, 32'h43238fde} /* (15, 0, 30) {real, imag} */,
  {32'hc1363970, 32'h42c3a941} /* (15, 0, 29) {real, imag} */,
  {32'hc1f757ba, 32'h42913e16} /* (15, 0, 28) {real, imag} */,
  {32'hc2df31fc, 32'hc14dea82} /* (15, 0, 27) {real, imag} */,
  {32'h4022ef10, 32'h4298c1df} /* (15, 0, 26) {real, imag} */,
  {32'hc28d10d7, 32'hc20e30e3} /* (15, 0, 25) {real, imag} */,
  {32'h420dc387, 32'hc219860f} /* (15, 0, 24) {real, imag} */,
  {32'hc2853214, 32'h417eefc4} /* (15, 0, 23) {real, imag} */,
  {32'hbe99e340, 32'hc2160fef} /* (15, 0, 22) {real, imag} */,
  {32'hc10fdaf2, 32'hc27b9c7e} /* (15, 0, 21) {real, imag} */,
  {32'hc229049c, 32'hc1f0c92e} /* (15, 0, 20) {real, imag} */,
  {32'h41158728, 32'hc17f065b} /* (15, 0, 19) {real, imag} */,
  {32'h41cb3ef5, 32'h4222f87b} /* (15, 0, 18) {real, imag} */,
  {32'h40cea744, 32'hc15d8c4e} /* (15, 0, 17) {real, imag} */,
  {32'h41832fd1, 32'h00000000} /* (15, 0, 16) {real, imag} */,
  {32'h40cea744, 32'h415d8c4e} /* (15, 0, 15) {real, imag} */,
  {32'h41cb3ef5, 32'hc222f87b} /* (15, 0, 14) {real, imag} */,
  {32'h41158728, 32'h417f065b} /* (15, 0, 13) {real, imag} */,
  {32'hc229049c, 32'h41f0c92e} /* (15, 0, 12) {real, imag} */,
  {32'hc10fdaf2, 32'h427b9c7e} /* (15, 0, 11) {real, imag} */,
  {32'hbe99e340, 32'h42160fef} /* (15, 0, 10) {real, imag} */,
  {32'hc2853214, 32'hc17eefc4} /* (15, 0, 9) {real, imag} */,
  {32'h420dc387, 32'h4219860f} /* (15, 0, 8) {real, imag} */,
  {32'hc28d10d7, 32'h420e30e3} /* (15, 0, 7) {real, imag} */,
  {32'h4022ef10, 32'hc298c1df} /* (15, 0, 6) {real, imag} */,
  {32'hc2df31fc, 32'h414dea82} /* (15, 0, 5) {real, imag} */,
  {32'hc1f757ba, 32'hc2913e16} /* (15, 0, 4) {real, imag} */,
  {32'hc1363970, 32'hc2c3a941} /* (15, 0, 3) {real, imag} */,
  {32'hc1f9e1d0, 32'hc3238fde} /* (15, 0, 2) {real, imag} */,
  {32'h4415afcb, 32'h442b896b} /* (15, 0, 1) {real, imag} */,
  {32'h443277c3, 32'h00000000} /* (15, 0, 0) {real, imag} */,
  {32'h44f3120e, 32'hc4a1e9ca} /* (14, 31, 31) {real, imag} */,
  {32'hc3e6e8f9, 32'h4390bc8c} /* (14, 31, 30) {real, imag} */,
  {32'hc19c3b90, 32'h42c3c85c} /* (14, 31, 29) {real, imag} */,
  {32'h42237202, 32'hc1c661b4} /* (14, 31, 28) {real, imag} */,
  {32'hc1ac1590, 32'h41585746} /* (14, 31, 27) {real, imag} */,
  {32'hc1c924a8, 32'h41d04472} /* (14, 31, 26) {real, imag} */,
  {32'hc08b2f70, 32'h42224089} /* (14, 31, 25) {real, imag} */,
  {32'h414c55b8, 32'h41a60edb} /* (14, 31, 24) {real, imag} */,
  {32'hc208378b, 32'h41c32a29} /* (14, 31, 23) {real, imag} */,
  {32'h3e8fcf80, 32'hc262eb90} /* (14, 31, 22) {real, imag} */,
  {32'hc232eb28, 32'h4161f31f} /* (14, 31, 21) {real, imag} */,
  {32'h41cd5c36, 32'hc146a7a8} /* (14, 31, 20) {real, imag} */,
  {32'h417765ed, 32'hc2794f6e} /* (14, 31, 19) {real, imag} */,
  {32'hc26dedfa, 32'h3f52ad30} /* (14, 31, 18) {real, imag} */,
  {32'hc1a0f109, 32'h420ea118} /* (14, 31, 17) {real, imag} */,
  {32'h42681c11, 32'h00000000} /* (14, 31, 16) {real, imag} */,
  {32'hc1a0f109, 32'hc20ea118} /* (14, 31, 15) {real, imag} */,
  {32'hc26dedfa, 32'hbf52ad30} /* (14, 31, 14) {real, imag} */,
  {32'h417765ed, 32'h42794f6e} /* (14, 31, 13) {real, imag} */,
  {32'h41cd5c36, 32'h4146a7a8} /* (14, 31, 12) {real, imag} */,
  {32'hc232eb28, 32'hc161f31f} /* (14, 31, 11) {real, imag} */,
  {32'h3e8fcf80, 32'h4262eb90} /* (14, 31, 10) {real, imag} */,
  {32'hc208378b, 32'hc1c32a29} /* (14, 31, 9) {real, imag} */,
  {32'h414c55b8, 32'hc1a60edb} /* (14, 31, 8) {real, imag} */,
  {32'hc08b2f70, 32'hc2224089} /* (14, 31, 7) {real, imag} */,
  {32'hc1c924a8, 32'hc1d04472} /* (14, 31, 6) {real, imag} */,
  {32'hc1ac1590, 32'hc1585746} /* (14, 31, 5) {real, imag} */,
  {32'h42237202, 32'h41c661b4} /* (14, 31, 4) {real, imag} */,
  {32'hc19c3b90, 32'hc2c3c85c} /* (14, 31, 3) {real, imag} */,
  {32'hc3e6e8f9, 32'hc390bc8c} /* (14, 31, 2) {real, imag} */,
  {32'h44f3120e, 32'h44a1e9ca} /* (14, 31, 1) {real, imag} */,
  {32'h451a6f8e, 32'h00000000} /* (14, 31, 0) {real, imag} */,
  {32'h45157487, 32'hc493bace} /* (14, 30, 31) {real, imag} */,
  {32'hc46858c5, 32'h4337a81f} /* (14, 30, 30) {real, imag} */,
  {32'h426c9417, 32'h4303f189} /* (14, 30, 29) {real, imag} */,
  {32'h434a2995, 32'h40e6df50} /* (14, 30, 28) {real, imag} */,
  {32'hc2081c6c, 32'h410d0d2a} /* (14, 30, 27) {real, imag} */,
  {32'h4227e94a, 32'hc2d9ebef} /* (14, 30, 26) {real, imag} */,
  {32'hc0db5be8, 32'h42831f14} /* (14, 30, 25) {real, imag} */,
  {32'h422c7be5, 32'h42b593ee} /* (14, 30, 24) {real, imag} */,
  {32'hc29dd30a, 32'hc11e4494} /* (14, 30, 23) {real, imag} */,
  {32'h43030f37, 32'h4289f147} /* (14, 30, 22) {real, imag} */,
  {32'hc068d368, 32'h42637e56} /* (14, 30, 21) {real, imag} */,
  {32'h428b9e29, 32'h406c4430} /* (14, 30, 20) {real, imag} */,
  {32'hc2675ba0, 32'hc2117978} /* (14, 30, 19) {real, imag} */,
  {32'h400eb058, 32'h425fc270} /* (14, 30, 18) {real, imag} */,
  {32'h41b9c76c, 32'h426a8110} /* (14, 30, 17) {real, imag} */,
  {32'h42450735, 32'h00000000} /* (14, 30, 16) {real, imag} */,
  {32'h41b9c76c, 32'hc26a8110} /* (14, 30, 15) {real, imag} */,
  {32'h400eb058, 32'hc25fc270} /* (14, 30, 14) {real, imag} */,
  {32'hc2675ba0, 32'h42117978} /* (14, 30, 13) {real, imag} */,
  {32'h428b9e29, 32'hc06c4430} /* (14, 30, 12) {real, imag} */,
  {32'hc068d368, 32'hc2637e56} /* (14, 30, 11) {real, imag} */,
  {32'h43030f37, 32'hc289f147} /* (14, 30, 10) {real, imag} */,
  {32'hc29dd30a, 32'h411e4494} /* (14, 30, 9) {real, imag} */,
  {32'h422c7be5, 32'hc2b593ee} /* (14, 30, 8) {real, imag} */,
  {32'hc0db5be8, 32'hc2831f14} /* (14, 30, 7) {real, imag} */,
  {32'h4227e94a, 32'h42d9ebef} /* (14, 30, 6) {real, imag} */,
  {32'hc2081c6c, 32'hc10d0d2a} /* (14, 30, 5) {real, imag} */,
  {32'h434a2995, 32'hc0e6df50} /* (14, 30, 4) {real, imag} */,
  {32'h426c9417, 32'hc303f189} /* (14, 30, 3) {real, imag} */,
  {32'hc46858c5, 32'hc337a81f} /* (14, 30, 2) {real, imag} */,
  {32'h45157487, 32'h4493bace} /* (14, 30, 1) {real, imag} */,
  {32'h451ebfd6, 32'h00000000} /* (14, 30, 0) {real, imag} */,
  {32'h451a9d66, 32'hc43ff838} /* (14, 29, 31) {real, imag} */,
  {32'hc45c8030, 32'h43109618} /* (14, 29, 30) {real, imag} */,
  {32'h427a3e93, 32'h428c97f8} /* (14, 29, 29) {real, imag} */,
  {32'h42aa35d8, 32'hc21efe4f} /* (14, 29, 28) {real, imag} */,
  {32'hc1c04220, 32'hc05c4cb0} /* (14, 29, 27) {real, imag} */,
  {32'h429c3d9a, 32'h40afbba2} /* (14, 29, 26) {real, imag} */,
  {32'h431b73bb, 32'h4284a81c} /* (14, 29, 25) {real, imag} */,
  {32'h40dac28a, 32'h42b5978d} /* (14, 29, 24) {real, imag} */,
  {32'hc24ec9ae, 32'h41fb5852} /* (14, 29, 23) {real, imag} */,
  {32'hc18c4af4, 32'h42e3f65c} /* (14, 29, 22) {real, imag} */,
  {32'hc20ab5d8, 32'h4246279d} /* (14, 29, 21) {real, imag} */,
  {32'h410694a8, 32'h4183d635} /* (14, 29, 20) {real, imag} */,
  {32'h4149e7c4, 32'h42b19d8a} /* (14, 29, 19) {real, imag} */,
  {32'hc0ff5c20, 32'h42b2cadd} /* (14, 29, 18) {real, imag} */,
  {32'h3c829000, 32'hc20d2efe} /* (14, 29, 17) {real, imag} */,
  {32'hc2b5a5f6, 32'h00000000} /* (14, 29, 16) {real, imag} */,
  {32'h3c829000, 32'h420d2efe} /* (14, 29, 15) {real, imag} */,
  {32'hc0ff5c20, 32'hc2b2cadd} /* (14, 29, 14) {real, imag} */,
  {32'h4149e7c4, 32'hc2b19d8a} /* (14, 29, 13) {real, imag} */,
  {32'h410694a8, 32'hc183d635} /* (14, 29, 12) {real, imag} */,
  {32'hc20ab5d8, 32'hc246279d} /* (14, 29, 11) {real, imag} */,
  {32'hc18c4af4, 32'hc2e3f65c} /* (14, 29, 10) {real, imag} */,
  {32'hc24ec9ae, 32'hc1fb5852} /* (14, 29, 9) {real, imag} */,
  {32'h40dac28a, 32'hc2b5978d} /* (14, 29, 8) {real, imag} */,
  {32'h431b73bb, 32'hc284a81c} /* (14, 29, 7) {real, imag} */,
  {32'h429c3d9a, 32'hc0afbba2} /* (14, 29, 6) {real, imag} */,
  {32'hc1c04220, 32'h405c4cb0} /* (14, 29, 5) {real, imag} */,
  {32'h42aa35d8, 32'h421efe4f} /* (14, 29, 4) {real, imag} */,
  {32'h427a3e93, 32'hc28c97f8} /* (14, 29, 3) {real, imag} */,
  {32'hc45c8030, 32'hc3109618} /* (14, 29, 2) {real, imag} */,
  {32'h451a9d66, 32'h443ff838} /* (14, 29, 1) {real, imag} */,
  {32'h452149c2, 32'h00000000} /* (14, 29, 0) {real, imag} */,
  {32'h45181b21, 32'hc411fa9b} /* (14, 28, 31) {real, imag} */,
  {32'hc4839fd8, 32'h42f5e508} /* (14, 28, 30) {real, imag} */,
  {32'h42b183bd, 32'hc227ed10} /* (14, 28, 29) {real, imag} */,
  {32'hc18657ac, 32'hc2faf042} /* (14, 28, 28) {real, imag} */,
  {32'hc24e8b36, 32'h431825a0} /* (14, 28, 27) {real, imag} */,
  {32'h40202460, 32'hc1b8453e} /* (14, 28, 26) {real, imag} */,
  {32'h42fc849b, 32'hbf918180} /* (14, 28, 25) {real, imag} */,
  {32'h3ff06758, 32'h4283eb76} /* (14, 28, 24) {real, imag} */,
  {32'hc2b06890, 32'h41b4bc44} /* (14, 28, 23) {real, imag} */,
  {32'hc14eece0, 32'hc2cd8d08} /* (14, 28, 22) {real, imag} */,
  {32'h423e1224, 32'h4264a7de} /* (14, 28, 21) {real, imag} */,
  {32'hc1d4a852, 32'h41e3ed07} /* (14, 28, 20) {real, imag} */,
  {32'h41bae2df, 32'hc159e710} /* (14, 28, 19) {real, imag} */,
  {32'hc1afddd4, 32'h421eb019} /* (14, 28, 18) {real, imag} */,
  {32'h4211e41f, 32'h4092c938} /* (14, 28, 17) {real, imag} */,
  {32'hc19f87c1, 32'h00000000} /* (14, 28, 16) {real, imag} */,
  {32'h4211e41f, 32'hc092c938} /* (14, 28, 15) {real, imag} */,
  {32'hc1afddd4, 32'hc21eb019} /* (14, 28, 14) {real, imag} */,
  {32'h41bae2df, 32'h4159e710} /* (14, 28, 13) {real, imag} */,
  {32'hc1d4a852, 32'hc1e3ed07} /* (14, 28, 12) {real, imag} */,
  {32'h423e1224, 32'hc264a7de} /* (14, 28, 11) {real, imag} */,
  {32'hc14eece0, 32'h42cd8d08} /* (14, 28, 10) {real, imag} */,
  {32'hc2b06890, 32'hc1b4bc44} /* (14, 28, 9) {real, imag} */,
  {32'h3ff06758, 32'hc283eb76} /* (14, 28, 8) {real, imag} */,
  {32'h42fc849b, 32'h3f918180} /* (14, 28, 7) {real, imag} */,
  {32'h40202460, 32'h41b8453e} /* (14, 28, 6) {real, imag} */,
  {32'hc24e8b36, 32'hc31825a0} /* (14, 28, 5) {real, imag} */,
  {32'hc18657ac, 32'h42faf042} /* (14, 28, 4) {real, imag} */,
  {32'h42b183bd, 32'h4227ed10} /* (14, 28, 3) {real, imag} */,
  {32'hc4839fd8, 32'hc2f5e508} /* (14, 28, 2) {real, imag} */,
  {32'h45181b21, 32'h4411fa9b} /* (14, 28, 1) {real, imag} */,
  {32'h4523b8b1, 32'h00000000} /* (14, 28, 0) {real, imag} */,
  {32'h4519c6cf, 32'hc41d6277} /* (14, 27, 31) {real, imag} */,
  {32'hc4887f53, 32'h43686a51} /* (14, 27, 30) {real, imag} */,
  {32'hc20255af, 32'hc3011b4c} /* (14, 27, 29) {real, imag} */,
  {32'h42795972, 32'hc3a38308} /* (14, 27, 28) {real, imag} */,
  {32'hc30d4274, 32'h433428b2} /* (14, 27, 27) {real, imag} */,
  {32'hc2aa4c00, 32'hbf8988a0} /* (14, 27, 26) {real, imag} */,
  {32'hc1744134, 32'hc255d29e} /* (14, 27, 25) {real, imag} */,
  {32'hc29e4f78, 32'h4340f148} /* (14, 27, 24) {real, imag} */,
  {32'hc2e827b5, 32'h40c2be64} /* (14, 27, 23) {real, imag} */,
  {32'h421153d7, 32'hc2fc2cfa} /* (14, 27, 22) {real, imag} */,
  {32'h41b5921f, 32'h430db24a} /* (14, 27, 21) {real, imag} */,
  {32'hc1ab20de, 32'hc26b03c8} /* (14, 27, 20) {real, imag} */,
  {32'h428ded5a, 32'hc22973b8} /* (14, 27, 19) {real, imag} */,
  {32'hc2aca7ed, 32'h424fe81e} /* (14, 27, 18) {real, imag} */,
  {32'h4251d5d9, 32'hc2049f3e} /* (14, 27, 17) {real, imag} */,
  {32'h42cb09b2, 32'h00000000} /* (14, 27, 16) {real, imag} */,
  {32'h4251d5d9, 32'h42049f3e} /* (14, 27, 15) {real, imag} */,
  {32'hc2aca7ed, 32'hc24fe81e} /* (14, 27, 14) {real, imag} */,
  {32'h428ded5a, 32'h422973b8} /* (14, 27, 13) {real, imag} */,
  {32'hc1ab20de, 32'h426b03c8} /* (14, 27, 12) {real, imag} */,
  {32'h41b5921f, 32'hc30db24a} /* (14, 27, 11) {real, imag} */,
  {32'h421153d7, 32'h42fc2cfa} /* (14, 27, 10) {real, imag} */,
  {32'hc2e827b5, 32'hc0c2be64} /* (14, 27, 9) {real, imag} */,
  {32'hc29e4f78, 32'hc340f148} /* (14, 27, 8) {real, imag} */,
  {32'hc1744134, 32'h4255d29e} /* (14, 27, 7) {real, imag} */,
  {32'hc2aa4c00, 32'h3f8988a0} /* (14, 27, 6) {real, imag} */,
  {32'hc30d4274, 32'hc33428b2} /* (14, 27, 5) {real, imag} */,
  {32'h42795972, 32'h43a38308} /* (14, 27, 4) {real, imag} */,
  {32'hc20255af, 32'h43011b4c} /* (14, 27, 3) {real, imag} */,
  {32'hc4887f53, 32'hc3686a51} /* (14, 27, 2) {real, imag} */,
  {32'h4519c6cf, 32'h441d6277} /* (14, 27, 1) {real, imag} */,
  {32'h45249dc7, 32'h00000000} /* (14, 27, 0) {real, imag} */,
  {32'h45229fee, 32'hc3eaa004} /* (14, 26, 31) {real, imag} */,
  {32'hc49036d2, 32'h43808881} /* (14, 26, 30) {real, imag} */,
  {32'hc2fc3c81, 32'hc2ab8fe4} /* (14, 26, 29) {real, imag} */,
  {32'h42208ee0, 32'hc30e861c} /* (14, 26, 28) {real, imag} */,
  {32'hc21805be, 32'h432d708f} /* (14, 26, 27) {real, imag} */,
  {32'hc22ee8cc, 32'h42d2ad62} /* (14, 26, 26) {real, imag} */,
  {32'hc238168e, 32'h4284b0b9} /* (14, 26, 25) {real, imag} */,
  {32'hc2304444, 32'h42414ca6} /* (14, 26, 24) {real, imag} */,
  {32'h43060d30, 32'hc248b4b2} /* (14, 26, 23) {real, imag} */,
  {32'h40a5f618, 32'hc29bb1b4} /* (14, 26, 22) {real, imag} */,
  {32'hc18cb7fe, 32'h4212f57e} /* (14, 26, 21) {real, imag} */,
  {32'hc20b4417, 32'h40effa20} /* (14, 26, 20) {real, imag} */,
  {32'h42d01edf, 32'hbfc571b0} /* (14, 26, 19) {real, imag} */,
  {32'hc27966c2, 32'h4238b0f3} /* (14, 26, 18) {real, imag} */,
  {32'h427ba604, 32'hc28365f0} /* (14, 26, 17) {real, imag} */,
  {32'hc08281c0, 32'h00000000} /* (14, 26, 16) {real, imag} */,
  {32'h427ba604, 32'h428365f0} /* (14, 26, 15) {real, imag} */,
  {32'hc27966c2, 32'hc238b0f3} /* (14, 26, 14) {real, imag} */,
  {32'h42d01edf, 32'h3fc571b0} /* (14, 26, 13) {real, imag} */,
  {32'hc20b4417, 32'hc0effa20} /* (14, 26, 12) {real, imag} */,
  {32'hc18cb7fe, 32'hc212f57e} /* (14, 26, 11) {real, imag} */,
  {32'h40a5f618, 32'h429bb1b4} /* (14, 26, 10) {real, imag} */,
  {32'h43060d30, 32'h4248b4b2} /* (14, 26, 9) {real, imag} */,
  {32'hc2304444, 32'hc2414ca6} /* (14, 26, 8) {real, imag} */,
  {32'hc238168e, 32'hc284b0b9} /* (14, 26, 7) {real, imag} */,
  {32'hc22ee8cc, 32'hc2d2ad62} /* (14, 26, 6) {real, imag} */,
  {32'hc21805be, 32'hc32d708f} /* (14, 26, 5) {real, imag} */,
  {32'h42208ee0, 32'h430e861c} /* (14, 26, 4) {real, imag} */,
  {32'hc2fc3c81, 32'h42ab8fe4} /* (14, 26, 3) {real, imag} */,
  {32'hc49036d2, 32'hc3808881} /* (14, 26, 2) {real, imag} */,
  {32'h45229fee, 32'h43eaa004} /* (14, 26, 1) {real, imag} */,
  {32'h451693d3, 32'h00000000} /* (14, 26, 0) {real, imag} */,
  {32'h45257c8b, 32'hc3f087fc} /* (14, 25, 31) {real, imag} */,
  {32'hc4984704, 32'h43682560} /* (14, 25, 30) {real, imag} */,
  {32'h41c6ec0a, 32'hc2283eb8} /* (14, 25, 29) {real, imag} */,
  {32'h42bf6a38, 32'hc2d60a41} /* (14, 25, 28) {real, imag} */,
  {32'hc3611ef6, 32'h42e88991} /* (14, 25, 27) {real, imag} */,
  {32'h4275da5a, 32'hc0054c10} /* (14, 25, 26) {real, imag} */,
  {32'h41a78410, 32'h42a31e89} /* (14, 25, 25) {real, imag} */,
  {32'hc2e25446, 32'h427e5442} /* (14, 25, 24) {real, imag} */,
  {32'h42a78ea1, 32'hc20d765e} /* (14, 25, 23) {real, imag} */,
  {32'hc2f89de0, 32'hc18fd3ca} /* (14, 25, 22) {real, imag} */,
  {32'hc215f34b, 32'h427750da} /* (14, 25, 21) {real, imag} */,
  {32'h40cce074, 32'h428fb8ec} /* (14, 25, 20) {real, imag} */,
  {32'h40159d68, 32'h42742eb3} /* (14, 25, 19) {real, imag} */,
  {32'h41d1daf6, 32'h407c9850} /* (14, 25, 18) {real, imag} */,
  {32'hc139dfe5, 32'h425f1efc} /* (14, 25, 17) {real, imag} */,
  {32'hc282a708, 32'h00000000} /* (14, 25, 16) {real, imag} */,
  {32'hc139dfe5, 32'hc25f1efc} /* (14, 25, 15) {real, imag} */,
  {32'h41d1daf6, 32'hc07c9850} /* (14, 25, 14) {real, imag} */,
  {32'h40159d68, 32'hc2742eb3} /* (14, 25, 13) {real, imag} */,
  {32'h40cce074, 32'hc28fb8ec} /* (14, 25, 12) {real, imag} */,
  {32'hc215f34b, 32'hc27750da} /* (14, 25, 11) {real, imag} */,
  {32'hc2f89de0, 32'h418fd3ca} /* (14, 25, 10) {real, imag} */,
  {32'h42a78ea1, 32'h420d765e} /* (14, 25, 9) {real, imag} */,
  {32'hc2e25446, 32'hc27e5442} /* (14, 25, 8) {real, imag} */,
  {32'h41a78410, 32'hc2a31e89} /* (14, 25, 7) {real, imag} */,
  {32'h4275da5a, 32'h40054c10} /* (14, 25, 6) {real, imag} */,
  {32'hc3611ef6, 32'hc2e88991} /* (14, 25, 5) {real, imag} */,
  {32'h42bf6a38, 32'h42d60a41} /* (14, 25, 4) {real, imag} */,
  {32'h41c6ec0a, 32'h42283eb8} /* (14, 25, 3) {real, imag} */,
  {32'hc4984704, 32'hc3682560} /* (14, 25, 2) {real, imag} */,
  {32'h45257c8b, 32'h43f087fc} /* (14, 25, 1) {real, imag} */,
  {32'h45063682, 32'h00000000} /* (14, 25, 0) {real, imag} */,
  {32'h4519b710, 32'hc3cf621a} /* (14, 24, 31) {real, imag} */,
  {32'hc4898d34, 32'h43ba2558} /* (14, 24, 30) {real, imag} */,
  {32'h41c46cde, 32'hc33b7c8f} /* (14, 24, 29) {real, imag} */,
  {32'h43222fde, 32'hc33f4b6b} /* (14, 24, 28) {real, imag} */,
  {32'hc3816bb6, 32'h43322795} /* (14, 24, 27) {real, imag} */,
  {32'hc30e5f6a, 32'h3fe89e00} /* (14, 24, 26) {real, imag} */,
  {32'h431bc801, 32'hc28576df} /* (14, 24, 25) {real, imag} */,
  {32'h4221ed74, 32'hc1ad5092} /* (14, 24, 24) {real, imag} */,
  {32'h42643858, 32'hc1af07e0} /* (14, 24, 23) {real, imag} */,
  {32'hc2521334, 32'hc2836a68} /* (14, 24, 22) {real, imag} */,
  {32'hc25624bc, 32'h420684ec} /* (14, 24, 21) {real, imag} */,
  {32'hc28774d2, 32'h42341d3e} /* (14, 24, 20) {real, imag} */,
  {32'hc2428e0c, 32'hbfd880f0} /* (14, 24, 19) {real, imag} */,
  {32'hc2ee75a9, 32'h409be9a0} /* (14, 24, 18) {real, imag} */,
  {32'hc2c1b31c, 32'h42777724} /* (14, 24, 17) {real, imag} */,
  {32'hc1718c32, 32'h00000000} /* (14, 24, 16) {real, imag} */,
  {32'hc2c1b31c, 32'hc2777724} /* (14, 24, 15) {real, imag} */,
  {32'hc2ee75a9, 32'hc09be9a0} /* (14, 24, 14) {real, imag} */,
  {32'hc2428e0c, 32'h3fd880f0} /* (14, 24, 13) {real, imag} */,
  {32'hc28774d2, 32'hc2341d3e} /* (14, 24, 12) {real, imag} */,
  {32'hc25624bc, 32'hc20684ec} /* (14, 24, 11) {real, imag} */,
  {32'hc2521334, 32'h42836a68} /* (14, 24, 10) {real, imag} */,
  {32'h42643858, 32'h41af07e0} /* (14, 24, 9) {real, imag} */,
  {32'h4221ed74, 32'h41ad5092} /* (14, 24, 8) {real, imag} */,
  {32'h431bc801, 32'h428576df} /* (14, 24, 7) {real, imag} */,
  {32'hc30e5f6a, 32'hbfe89e00} /* (14, 24, 6) {real, imag} */,
  {32'hc3816bb6, 32'hc3322795} /* (14, 24, 5) {real, imag} */,
  {32'h43222fde, 32'h433f4b6b} /* (14, 24, 4) {real, imag} */,
  {32'h41c46cde, 32'h433b7c8f} /* (14, 24, 3) {real, imag} */,
  {32'hc4898d34, 32'hc3ba2558} /* (14, 24, 2) {real, imag} */,
  {32'h4519b710, 32'h43cf621a} /* (14, 24, 1) {real, imag} */,
  {32'h44e49fb3, 32'h00000000} /* (14, 24, 0) {real, imag} */,
  {32'h44fe9254, 32'hc388e780} /* (14, 23, 31) {real, imag} */,
  {32'hc467c811, 32'h4373f35c} /* (14, 23, 30) {real, imag} */,
  {32'h426d37a9, 32'hc326bfc2} /* (14, 23, 29) {real, imag} */,
  {32'h4303c72e, 32'hc3249cd6} /* (14, 23, 28) {real, imag} */,
  {32'hc3352074, 32'h42952570} /* (14, 23, 27) {real, imag} */,
  {32'hc0fb8580, 32'hc14d421a} /* (14, 23, 26) {real, imag} */,
  {32'h42fdd4f1, 32'h41dda000} /* (14, 23, 25) {real, imag} */,
  {32'hc20aebc5, 32'h4191762a} /* (14, 23, 24) {real, imag} */,
  {32'hc11c1d80, 32'h42e64c16} /* (14, 23, 23) {real, imag} */,
  {32'hc1f876a4, 32'hc2db8856} /* (14, 23, 22) {real, imag} */,
  {32'h424d8cee, 32'hc20e0b06} /* (14, 23, 21) {real, imag} */,
  {32'h42105eac, 32'h42107313} /* (14, 23, 20) {real, imag} */,
  {32'h41496bc2, 32'h423eb35a} /* (14, 23, 19) {real, imag} */,
  {32'hbfc36e68, 32'h428aa58f} /* (14, 23, 18) {real, imag} */,
  {32'h423a87b2, 32'h42213bd6} /* (14, 23, 17) {real, imag} */,
  {32'hc149cc16, 32'h00000000} /* (14, 23, 16) {real, imag} */,
  {32'h423a87b2, 32'hc2213bd6} /* (14, 23, 15) {real, imag} */,
  {32'hbfc36e68, 32'hc28aa58f} /* (14, 23, 14) {real, imag} */,
  {32'h41496bc2, 32'hc23eb35a} /* (14, 23, 13) {real, imag} */,
  {32'h42105eac, 32'hc2107313} /* (14, 23, 12) {real, imag} */,
  {32'h424d8cee, 32'h420e0b06} /* (14, 23, 11) {real, imag} */,
  {32'hc1f876a4, 32'h42db8856} /* (14, 23, 10) {real, imag} */,
  {32'hc11c1d80, 32'hc2e64c16} /* (14, 23, 9) {real, imag} */,
  {32'hc20aebc5, 32'hc191762a} /* (14, 23, 8) {real, imag} */,
  {32'h42fdd4f1, 32'hc1dda000} /* (14, 23, 7) {real, imag} */,
  {32'hc0fb8580, 32'h414d421a} /* (14, 23, 6) {real, imag} */,
  {32'hc3352074, 32'hc2952570} /* (14, 23, 5) {real, imag} */,
  {32'h4303c72e, 32'h43249cd6} /* (14, 23, 4) {real, imag} */,
  {32'h426d37a9, 32'h4326bfc2} /* (14, 23, 3) {real, imag} */,
  {32'hc467c811, 32'hc373f35c} /* (14, 23, 2) {real, imag} */,
  {32'h44fe9254, 32'h4388e780} /* (14, 23, 1) {real, imag} */,
  {32'h44aa08e2, 32'h00000000} /* (14, 23, 0) {real, imag} */,
  {32'h44b4b1a7, 32'hc3300817} /* (14, 22, 31) {real, imag} */,
  {32'hc421733d, 32'h432ab9d6} /* (14, 22, 30) {real, imag} */,
  {32'h413a4670, 32'hc32d93a4} /* (14, 22, 29) {real, imag} */,
  {32'h43159aa6, 32'hc365557e} /* (14, 22, 28) {real, imag} */,
  {32'hc33e53a0, 32'h42cb2c7a} /* (14, 22, 27) {real, imag} */,
  {32'hc28efbd0, 32'h42809522} /* (14, 22, 26) {real, imag} */,
  {32'h42f92e79, 32'h41ce29c9} /* (14, 22, 25) {real, imag} */,
  {32'hc2237ddc, 32'h42b5ed98} /* (14, 22, 24) {real, imag} */,
  {32'hc2d127de, 32'h43186f21} /* (14, 22, 23) {real, imag} */,
  {32'hc21cd015, 32'h421876ae} /* (14, 22, 22) {real, imag} */,
  {32'hc2d7be15, 32'hc2a1f628} /* (14, 22, 21) {real, imag} */,
  {32'h428259da, 32'hc29c7d36} /* (14, 22, 20) {real, imag} */,
  {32'h41d7db8f, 32'hc0bfd830} /* (14, 22, 19) {real, imag} */,
  {32'hc226cd0e, 32'h42438c8c} /* (14, 22, 18) {real, imag} */,
  {32'hc1b46e6a, 32'hc2e52132} /* (14, 22, 17) {real, imag} */,
  {32'h42804c96, 32'h00000000} /* (14, 22, 16) {real, imag} */,
  {32'hc1b46e6a, 32'h42e52132} /* (14, 22, 15) {real, imag} */,
  {32'hc226cd0e, 32'hc2438c8c} /* (14, 22, 14) {real, imag} */,
  {32'h41d7db8f, 32'h40bfd830} /* (14, 22, 13) {real, imag} */,
  {32'h428259da, 32'h429c7d36} /* (14, 22, 12) {real, imag} */,
  {32'hc2d7be15, 32'h42a1f628} /* (14, 22, 11) {real, imag} */,
  {32'hc21cd015, 32'hc21876ae} /* (14, 22, 10) {real, imag} */,
  {32'hc2d127de, 32'hc3186f21} /* (14, 22, 9) {real, imag} */,
  {32'hc2237ddc, 32'hc2b5ed98} /* (14, 22, 8) {real, imag} */,
  {32'h42f92e79, 32'hc1ce29c9} /* (14, 22, 7) {real, imag} */,
  {32'hc28efbd0, 32'hc2809522} /* (14, 22, 6) {real, imag} */,
  {32'hc33e53a0, 32'hc2cb2c7a} /* (14, 22, 5) {real, imag} */,
  {32'h43159aa6, 32'h4365557e} /* (14, 22, 4) {real, imag} */,
  {32'h413a4670, 32'h432d93a4} /* (14, 22, 3) {real, imag} */,
  {32'hc421733d, 32'hc32ab9d6} /* (14, 22, 2) {real, imag} */,
  {32'h44b4b1a7, 32'h43300817} /* (14, 22, 1) {real, imag} */,
  {32'h44983438, 32'h00000000} /* (14, 22, 0) {real, imag} */,
  {32'h43c06862, 32'h42a054c0} /* (14, 21, 31) {real, imag} */,
  {32'hc34af16d, 32'h4322a25f} /* (14, 21, 30) {real, imag} */,
  {32'h42ec9d13, 32'hc2f0fef9} /* (14, 21, 29) {real, imag} */,
  {32'h42ff8134, 32'hc2fdd604} /* (14, 21, 28) {real, imag} */,
  {32'hc3085644, 32'h42c35fe7} /* (14, 21, 27) {real, imag} */,
  {32'hc2cc8c9c, 32'h40354378} /* (14, 21, 26) {real, imag} */,
  {32'h41b46217, 32'hc2e2926d} /* (14, 21, 25) {real, imag} */,
  {32'h429206b5, 32'hc1b956c3} /* (14, 21, 24) {real, imag} */,
  {32'hbf83c7e0, 32'h424db68a} /* (14, 21, 23) {real, imag} */,
  {32'h412de2c8, 32'hc230d216} /* (14, 21, 22) {real, imag} */,
  {32'hc13fbb4c, 32'h40ea3cc4} /* (14, 21, 21) {real, imag} */,
  {32'hc135954b, 32'h430a888e} /* (14, 21, 20) {real, imag} */,
  {32'h420315d6, 32'h406a33a8} /* (14, 21, 19) {real, imag} */,
  {32'hc2884641, 32'hc25e1aac} /* (14, 21, 18) {real, imag} */,
  {32'hc204071a, 32'h417a60d4} /* (14, 21, 17) {real, imag} */,
  {32'hc22eb2b1, 32'h00000000} /* (14, 21, 16) {real, imag} */,
  {32'hc204071a, 32'hc17a60d4} /* (14, 21, 15) {real, imag} */,
  {32'hc2884641, 32'h425e1aac} /* (14, 21, 14) {real, imag} */,
  {32'h420315d6, 32'hc06a33a8} /* (14, 21, 13) {real, imag} */,
  {32'hc135954b, 32'hc30a888e} /* (14, 21, 12) {real, imag} */,
  {32'hc13fbb4c, 32'hc0ea3cc4} /* (14, 21, 11) {real, imag} */,
  {32'h412de2c8, 32'h4230d216} /* (14, 21, 10) {real, imag} */,
  {32'hbf83c7e0, 32'hc24db68a} /* (14, 21, 9) {real, imag} */,
  {32'h429206b5, 32'h41b956c3} /* (14, 21, 8) {real, imag} */,
  {32'h41b46217, 32'h42e2926d} /* (14, 21, 7) {real, imag} */,
  {32'hc2cc8c9c, 32'hc0354378} /* (14, 21, 6) {real, imag} */,
  {32'hc3085644, 32'hc2c35fe7} /* (14, 21, 5) {real, imag} */,
  {32'h42ff8134, 32'h42fdd604} /* (14, 21, 4) {real, imag} */,
  {32'h42ec9d13, 32'h42f0fef9} /* (14, 21, 3) {real, imag} */,
  {32'hc34af16d, 32'hc322a25f} /* (14, 21, 2) {real, imag} */,
  {32'h43c06862, 32'hc2a054c0} /* (14, 21, 1) {real, imag} */,
  {32'h44152456, 32'h00000000} /* (14, 21, 0) {real, imag} */,
  {32'hc47477ed, 32'h43674b40} /* (14, 20, 31) {real, imag} */,
  {32'h43ddeb3e, 32'h4141e300} /* (14, 20, 30) {real, imag} */,
  {32'h42f8d476, 32'hc1020434} /* (14, 20, 29) {real, imag} */,
  {32'hc0f606f0, 32'hc20ebf04} /* (14, 20, 28) {real, imag} */,
  {32'h41e55b10, 32'hc3067566} /* (14, 20, 27) {real, imag} */,
  {32'h420b2d90, 32'hc2fbf2c5} /* (14, 20, 26) {real, imag} */,
  {32'hc0cd1ad8, 32'hc218eacf} /* (14, 20, 25) {real, imag} */,
  {32'h421cfb38, 32'hc2901da6} /* (14, 20, 24) {real, imag} */,
  {32'hc29bf326, 32'hc03492cc} /* (14, 20, 23) {real, imag} */,
  {32'hc2d5bb9f, 32'h42bc5f00} /* (14, 20, 22) {real, imag} */,
  {32'h42bb628d, 32'h4213d66e} /* (14, 20, 21) {real, imag} */,
  {32'h42987bec, 32'h429a16df} /* (14, 20, 20) {real, imag} */,
  {32'hc2aef105, 32'h422df589} /* (14, 20, 19) {real, imag} */,
  {32'h4281b9da, 32'hc2e5cf5c} /* (14, 20, 18) {real, imag} */,
  {32'hc191a1ca, 32'h427c0db4} /* (14, 20, 17) {real, imag} */,
  {32'hc221fee5, 32'h00000000} /* (14, 20, 16) {real, imag} */,
  {32'hc191a1ca, 32'hc27c0db4} /* (14, 20, 15) {real, imag} */,
  {32'h4281b9da, 32'h42e5cf5c} /* (14, 20, 14) {real, imag} */,
  {32'hc2aef105, 32'hc22df589} /* (14, 20, 13) {real, imag} */,
  {32'h42987bec, 32'hc29a16df} /* (14, 20, 12) {real, imag} */,
  {32'h42bb628d, 32'hc213d66e} /* (14, 20, 11) {real, imag} */,
  {32'hc2d5bb9f, 32'hc2bc5f00} /* (14, 20, 10) {real, imag} */,
  {32'hc29bf326, 32'h403492cc} /* (14, 20, 9) {real, imag} */,
  {32'h421cfb38, 32'h42901da6} /* (14, 20, 8) {real, imag} */,
  {32'hc0cd1ad8, 32'h4218eacf} /* (14, 20, 7) {real, imag} */,
  {32'h420b2d90, 32'h42fbf2c5} /* (14, 20, 6) {real, imag} */,
  {32'h41e55b10, 32'h43067566} /* (14, 20, 5) {real, imag} */,
  {32'hc0f606f0, 32'h420ebf04} /* (14, 20, 4) {real, imag} */,
  {32'h42f8d476, 32'h41020434} /* (14, 20, 3) {real, imag} */,
  {32'h43ddeb3e, 32'hc141e300} /* (14, 20, 2) {real, imag} */,
  {32'hc47477ed, 32'hc3674b40} /* (14, 20, 1) {real, imag} */,
  {32'hc41197b0, 32'h00000000} /* (14, 20, 0) {real, imag} */,
  {32'hc4c6b476, 32'h4386b0c7} /* (14, 19, 31) {real, imag} */,
  {32'h4442fd8a, 32'hc2e0645a} /* (14, 19, 30) {real, imag} */,
  {32'h4362faab, 32'h4138ac20} /* (14, 19, 29) {real, imag} */,
  {32'hc3171922, 32'h429565ef} /* (14, 19, 28) {real, imag} */,
  {32'h42e2d35b, 32'hc310b76c} /* (14, 19, 27) {real, imag} */,
  {32'hc2a60bb6, 32'hc229b170} /* (14, 19, 26) {real, imag} */,
  {32'hc18bc170, 32'h42ae58cc} /* (14, 19, 25) {real, imag} */,
  {32'h42cacbcf, 32'h42431044} /* (14, 19, 24) {real, imag} */,
  {32'hc1b7b0b2, 32'h42150708} /* (14, 19, 23) {real, imag} */,
  {32'hc2adfd48, 32'hc29936a8} /* (14, 19, 22) {real, imag} */,
  {32'h42017e38, 32'hc2a8767b} /* (14, 19, 21) {real, imag} */,
  {32'h417eeb72, 32'hc1a8eb22} /* (14, 19, 20) {real, imag} */,
  {32'hc263e32e, 32'h4296dcc0} /* (14, 19, 19) {real, imag} */,
  {32'hc0eb6e10, 32'h41f6e2ec} /* (14, 19, 18) {real, imag} */,
  {32'h41154c40, 32'hc248dd78} /* (14, 19, 17) {real, imag} */,
  {32'h40522b00, 32'h00000000} /* (14, 19, 16) {real, imag} */,
  {32'h41154c40, 32'h4248dd78} /* (14, 19, 15) {real, imag} */,
  {32'hc0eb6e10, 32'hc1f6e2ec} /* (14, 19, 14) {real, imag} */,
  {32'hc263e32e, 32'hc296dcc0} /* (14, 19, 13) {real, imag} */,
  {32'h417eeb72, 32'h41a8eb22} /* (14, 19, 12) {real, imag} */,
  {32'h42017e38, 32'h42a8767b} /* (14, 19, 11) {real, imag} */,
  {32'hc2adfd48, 32'h429936a8} /* (14, 19, 10) {real, imag} */,
  {32'hc1b7b0b2, 32'hc2150708} /* (14, 19, 9) {real, imag} */,
  {32'h42cacbcf, 32'hc2431044} /* (14, 19, 8) {real, imag} */,
  {32'hc18bc170, 32'hc2ae58cc} /* (14, 19, 7) {real, imag} */,
  {32'hc2a60bb6, 32'h4229b170} /* (14, 19, 6) {real, imag} */,
  {32'h42e2d35b, 32'h4310b76c} /* (14, 19, 5) {real, imag} */,
  {32'hc3171922, 32'hc29565ef} /* (14, 19, 4) {real, imag} */,
  {32'h4362faab, 32'hc138ac20} /* (14, 19, 3) {real, imag} */,
  {32'h4442fd8a, 32'h42e0645a} /* (14, 19, 2) {real, imag} */,
  {32'hc4c6b476, 32'hc386b0c7} /* (14, 19, 1) {real, imag} */,
  {32'hc475c510, 32'h00000000} /* (14, 19, 0) {real, imag} */,
  {32'hc4f6d3dc, 32'h43921bed} /* (14, 18, 31) {real, imag} */,
  {32'h4455d7f0, 32'hc381e218} /* (14, 18, 30) {real, imag} */,
  {32'h4308cccc, 32'hc26c5253} /* (14, 18, 29) {real, imag} */,
  {32'hc311d9f3, 32'h43025cd5} /* (14, 18, 28) {real, imag} */,
  {32'h425e36ee, 32'hc181602e} /* (14, 18, 27) {real, imag} */,
  {32'hc2a35503, 32'hc207bcee} /* (14, 18, 26) {real, imag} */,
  {32'hc2e38beb, 32'h41f82068} /* (14, 18, 25) {real, imag} */,
  {32'h4252a9d9, 32'hc21ca296} /* (14, 18, 24) {real, imag} */,
  {32'hc208dca2, 32'hc1d338c4} /* (14, 18, 23) {real, imag} */,
  {32'h412af075, 32'hc247f048} /* (14, 18, 22) {real, imag} */,
  {32'hc2cb8484, 32'hc28aec35} /* (14, 18, 21) {real, imag} */,
  {32'h42248e3a, 32'hc26340bd} /* (14, 18, 20) {real, imag} */,
  {32'h41bdb0ee, 32'hc20f5cba} /* (14, 18, 19) {real, imag} */,
  {32'h42c5ff14, 32'hc2a2a4d1} /* (14, 18, 18) {real, imag} */,
  {32'h42b14f5d, 32'h4089d500} /* (14, 18, 17) {real, imag} */,
  {32'h40ff6460, 32'h00000000} /* (14, 18, 16) {real, imag} */,
  {32'h42b14f5d, 32'hc089d500} /* (14, 18, 15) {real, imag} */,
  {32'h42c5ff14, 32'h42a2a4d1} /* (14, 18, 14) {real, imag} */,
  {32'h41bdb0ee, 32'h420f5cba} /* (14, 18, 13) {real, imag} */,
  {32'h42248e3a, 32'h426340bd} /* (14, 18, 12) {real, imag} */,
  {32'hc2cb8484, 32'h428aec35} /* (14, 18, 11) {real, imag} */,
  {32'h412af075, 32'h4247f048} /* (14, 18, 10) {real, imag} */,
  {32'hc208dca2, 32'h41d338c4} /* (14, 18, 9) {real, imag} */,
  {32'h4252a9d9, 32'h421ca296} /* (14, 18, 8) {real, imag} */,
  {32'hc2e38beb, 32'hc1f82068} /* (14, 18, 7) {real, imag} */,
  {32'hc2a35503, 32'h4207bcee} /* (14, 18, 6) {real, imag} */,
  {32'h425e36ee, 32'h4181602e} /* (14, 18, 5) {real, imag} */,
  {32'hc311d9f3, 32'hc3025cd5} /* (14, 18, 4) {real, imag} */,
  {32'h4308cccc, 32'h426c5253} /* (14, 18, 3) {real, imag} */,
  {32'h4455d7f0, 32'h4381e218} /* (14, 18, 2) {real, imag} */,
  {32'hc4f6d3dc, 32'hc3921bed} /* (14, 18, 1) {real, imag} */,
  {32'hc4a6ce38, 32'h00000000} /* (14, 18, 0) {real, imag} */,
  {32'hc50b6eb6, 32'h435a8902} /* (14, 17, 31) {real, imag} */,
  {32'h4483c118, 32'hc34f7e2a} /* (14, 17, 30) {real, imag} */,
  {32'h4311d72d, 32'hc320246b} /* (14, 17, 29) {real, imag} */,
  {32'hc318e79c, 32'h4318d274} /* (14, 17, 28) {real, imag} */,
  {32'h42f69eb2, 32'h4182c4f5} /* (14, 17, 27) {real, imag} */,
  {32'hc3550d82, 32'hc1fa8060} /* (14, 17, 26) {real, imag} */,
  {32'hc2917e57, 32'hc2651a2a} /* (14, 17, 25) {real, imag} */,
  {32'h42d880e9, 32'hc2dbe528} /* (14, 17, 24) {real, imag} */,
  {32'h40ffdec0, 32'hc1d15d6f} /* (14, 17, 23) {real, imag} */,
  {32'h42655940, 32'hc2064c16} /* (14, 17, 22) {real, imag} */,
  {32'h42031f65, 32'hc0c64230} /* (14, 17, 21) {real, imag} */,
  {32'h41efe528, 32'hc2371ff1} /* (14, 17, 20) {real, imag} */,
  {32'hc28539d2, 32'hc254be30} /* (14, 17, 19) {real, imag} */,
  {32'hc1db872a, 32'hc06c0aa4} /* (14, 17, 18) {real, imag} */,
  {32'hc10fb39a, 32'h42922c44} /* (14, 17, 17) {real, imag} */,
  {32'h42279b7c, 32'h00000000} /* (14, 17, 16) {real, imag} */,
  {32'hc10fb39a, 32'hc2922c44} /* (14, 17, 15) {real, imag} */,
  {32'hc1db872a, 32'h406c0aa4} /* (14, 17, 14) {real, imag} */,
  {32'hc28539d2, 32'h4254be30} /* (14, 17, 13) {real, imag} */,
  {32'h41efe528, 32'h42371ff1} /* (14, 17, 12) {real, imag} */,
  {32'h42031f65, 32'h40c64230} /* (14, 17, 11) {real, imag} */,
  {32'h42655940, 32'h42064c16} /* (14, 17, 10) {real, imag} */,
  {32'h40ffdec0, 32'h41d15d6f} /* (14, 17, 9) {real, imag} */,
  {32'h42d880e9, 32'h42dbe528} /* (14, 17, 8) {real, imag} */,
  {32'hc2917e57, 32'h42651a2a} /* (14, 17, 7) {real, imag} */,
  {32'hc3550d82, 32'h41fa8060} /* (14, 17, 6) {real, imag} */,
  {32'h42f69eb2, 32'hc182c4f5} /* (14, 17, 5) {real, imag} */,
  {32'hc318e79c, 32'hc318d274} /* (14, 17, 4) {real, imag} */,
  {32'h4311d72d, 32'h4320246b} /* (14, 17, 3) {real, imag} */,
  {32'h4483c118, 32'h434f7e2a} /* (14, 17, 2) {real, imag} */,
  {32'hc50b6eb6, 32'hc35a8902} /* (14, 17, 1) {real, imag} */,
  {32'hc4e53322, 32'h00000000} /* (14, 17, 0) {real, imag} */,
  {32'hc51badd4, 32'h43c0a560} /* (14, 16, 31) {real, imag} */,
  {32'h448dfabd, 32'hc386087f} /* (14, 16, 30) {real, imag} */,
  {32'h42932dca, 32'hc32e91c5} /* (14, 16, 29) {real, imag} */,
  {32'hc31528a2, 32'h438e612c} /* (14, 16, 28) {real, imag} */,
  {32'h431ce952, 32'hc2ae9e2c} /* (14, 16, 27) {real, imag} */,
  {32'h41da6c7a, 32'hc2891eec} /* (14, 16, 26) {real, imag} */,
  {32'hc281ebf7, 32'h4187d08c} /* (14, 16, 25) {real, imag} */,
  {32'h42859c07, 32'h4279fd17} /* (14, 16, 24) {real, imag} */,
  {32'h42464378, 32'hc213c785} /* (14, 16, 23) {real, imag} */,
  {32'hbf51ab38, 32'hc2774f2e} /* (14, 16, 22) {real, imag} */,
  {32'h42a46a18, 32'hc2b8aebc} /* (14, 16, 21) {real, imag} */,
  {32'hc14049d5, 32'h42c0102e} /* (14, 16, 20) {real, imag} */,
  {32'hc2b2b8aa, 32'h429abefd} /* (14, 16, 19) {real, imag} */,
  {32'h4105702a, 32'h41a36260} /* (14, 16, 18) {real, imag} */,
  {32'h4082c780, 32'h41ac232e} /* (14, 16, 17) {real, imag} */,
  {32'hc14fa25c, 32'h00000000} /* (14, 16, 16) {real, imag} */,
  {32'h4082c780, 32'hc1ac232e} /* (14, 16, 15) {real, imag} */,
  {32'h4105702a, 32'hc1a36260} /* (14, 16, 14) {real, imag} */,
  {32'hc2b2b8aa, 32'hc29abefd} /* (14, 16, 13) {real, imag} */,
  {32'hc14049d5, 32'hc2c0102e} /* (14, 16, 12) {real, imag} */,
  {32'h42a46a18, 32'h42b8aebc} /* (14, 16, 11) {real, imag} */,
  {32'hbf51ab38, 32'h42774f2e} /* (14, 16, 10) {real, imag} */,
  {32'h42464378, 32'h4213c785} /* (14, 16, 9) {real, imag} */,
  {32'h42859c07, 32'hc279fd17} /* (14, 16, 8) {real, imag} */,
  {32'hc281ebf7, 32'hc187d08c} /* (14, 16, 7) {real, imag} */,
  {32'h41da6c7a, 32'h42891eec} /* (14, 16, 6) {real, imag} */,
  {32'h431ce952, 32'h42ae9e2c} /* (14, 16, 5) {real, imag} */,
  {32'hc31528a2, 32'hc38e612c} /* (14, 16, 4) {real, imag} */,
  {32'h42932dca, 32'h432e91c5} /* (14, 16, 3) {real, imag} */,
  {32'h448dfabd, 32'h4386087f} /* (14, 16, 2) {real, imag} */,
  {32'hc51badd4, 32'hc3c0a560} /* (14, 16, 1) {real, imag} */,
  {32'hc4db99c9, 32'h00000000} /* (14, 16, 0) {real, imag} */,
  {32'hc5249cee, 32'h43f758f3} /* (14, 15, 31) {real, imag} */,
  {32'h4487af84, 32'hc3697dae} /* (14, 15, 30) {real, imag} */,
  {32'h429035da, 32'hc2bffce6} /* (14, 15, 29) {real, imag} */,
  {32'hc30995f8, 32'h43935d28} /* (14, 15, 28) {real, imag} */,
  {32'h428f1cb2, 32'hc270318c} /* (14, 15, 27) {real, imag} */,
  {32'h41b87100, 32'hc389f6be} /* (14, 15, 26) {real, imag} */,
  {32'hc298e41f, 32'h42344c92} /* (14, 15, 25) {real, imag} */,
  {32'h434997a4, 32'hc1ec7738} /* (14, 15, 24) {real, imag} */,
  {32'h43027f5b, 32'hc22e7e80} /* (14, 15, 23) {real, imag} */,
  {32'hc28b8535, 32'hc2406f12} /* (14, 15, 22) {real, imag} */,
  {32'hc2a69dc0, 32'h42934561} /* (14, 15, 21) {real, imag} */,
  {32'h42256170, 32'h42888ca2} /* (14, 15, 20) {real, imag} */,
  {32'hc2e5e440, 32'hc2e8195c} /* (14, 15, 19) {real, imag} */,
  {32'hc21a1b0f, 32'hc150d3e9} /* (14, 15, 18) {real, imag} */,
  {32'hc22b7dfa, 32'h41b793a8} /* (14, 15, 17) {real, imag} */,
  {32'hc20ec7dc, 32'h00000000} /* (14, 15, 16) {real, imag} */,
  {32'hc22b7dfa, 32'hc1b793a8} /* (14, 15, 15) {real, imag} */,
  {32'hc21a1b0f, 32'h4150d3e9} /* (14, 15, 14) {real, imag} */,
  {32'hc2e5e440, 32'h42e8195c} /* (14, 15, 13) {real, imag} */,
  {32'h42256170, 32'hc2888ca2} /* (14, 15, 12) {real, imag} */,
  {32'hc2a69dc0, 32'hc2934561} /* (14, 15, 11) {real, imag} */,
  {32'hc28b8535, 32'h42406f12} /* (14, 15, 10) {real, imag} */,
  {32'h43027f5b, 32'h422e7e80} /* (14, 15, 9) {real, imag} */,
  {32'h434997a4, 32'h41ec7738} /* (14, 15, 8) {real, imag} */,
  {32'hc298e41f, 32'hc2344c92} /* (14, 15, 7) {real, imag} */,
  {32'h41b87100, 32'h4389f6be} /* (14, 15, 6) {real, imag} */,
  {32'h428f1cb2, 32'h4270318c} /* (14, 15, 5) {real, imag} */,
  {32'hc30995f8, 32'hc3935d28} /* (14, 15, 4) {real, imag} */,
  {32'h429035da, 32'h42bffce6} /* (14, 15, 3) {real, imag} */,
  {32'h4487af84, 32'h43697dae} /* (14, 15, 2) {real, imag} */,
  {32'hc5249cee, 32'hc3f758f3} /* (14, 15, 1) {real, imag} */,
  {32'hc4ed1ec4, 32'h00000000} /* (14, 15, 0) {real, imag} */,
  {32'hc520b3cc, 32'h43c886ff} /* (14, 14, 31) {real, imag} */,
  {32'h4457b00e, 32'hc3356b77} /* (14, 14, 30) {real, imag} */,
  {32'h4271a97e, 32'h41d29922} /* (14, 14, 29) {real, imag} */,
  {32'hc0cdde60, 32'h433aa18f} /* (14, 14, 28) {real, imag} */,
  {32'h431b1020, 32'hc2c0ebbc} /* (14, 14, 27) {real, imag} */,
  {32'h41fac247, 32'hc2d02ab9} /* (14, 14, 26) {real, imag} */,
  {32'hc2bad88d, 32'hc199b2d8} /* (14, 14, 25) {real, imag} */,
  {32'h42fe50d2, 32'h418430eb} /* (14, 14, 24) {real, imag} */,
  {32'h4162be36, 32'h3e42c400} /* (14, 14, 23) {real, imag} */,
  {32'hc1cbb10a, 32'h40c77564} /* (14, 14, 22) {real, imag} */,
  {32'hc1271d64, 32'hc2c32775} /* (14, 14, 21) {real, imag} */,
  {32'h4125e482, 32'hc1f95e42} /* (14, 14, 20) {real, imag} */,
  {32'hc108cbdc, 32'h422e9206} /* (14, 14, 19) {real, imag} */,
  {32'h411d4fcc, 32'hc105bab8} /* (14, 14, 18) {real, imag} */,
  {32'h427addde, 32'h428ec286} /* (14, 14, 17) {real, imag} */,
  {32'h4182cd1e, 32'h00000000} /* (14, 14, 16) {real, imag} */,
  {32'h427addde, 32'hc28ec286} /* (14, 14, 15) {real, imag} */,
  {32'h411d4fcc, 32'h4105bab8} /* (14, 14, 14) {real, imag} */,
  {32'hc108cbdc, 32'hc22e9206} /* (14, 14, 13) {real, imag} */,
  {32'h4125e482, 32'h41f95e42} /* (14, 14, 12) {real, imag} */,
  {32'hc1271d64, 32'h42c32775} /* (14, 14, 11) {real, imag} */,
  {32'hc1cbb10a, 32'hc0c77564} /* (14, 14, 10) {real, imag} */,
  {32'h4162be36, 32'hbe42c400} /* (14, 14, 9) {real, imag} */,
  {32'h42fe50d2, 32'hc18430eb} /* (14, 14, 8) {real, imag} */,
  {32'hc2bad88d, 32'h4199b2d8} /* (14, 14, 7) {real, imag} */,
  {32'h41fac247, 32'h42d02ab9} /* (14, 14, 6) {real, imag} */,
  {32'h431b1020, 32'h42c0ebbc} /* (14, 14, 5) {real, imag} */,
  {32'hc0cdde60, 32'hc33aa18f} /* (14, 14, 4) {real, imag} */,
  {32'h4271a97e, 32'hc1d29922} /* (14, 14, 3) {real, imag} */,
  {32'h4457b00e, 32'h43356b77} /* (14, 14, 2) {real, imag} */,
  {32'hc520b3cc, 32'hc3c886ff} /* (14, 14, 1) {real, imag} */,
  {32'hc4c9ba90, 32'h00000000} /* (14, 14, 0) {real, imag} */,
  {32'hc50c7100, 32'h4356be92} /* (14, 13, 31) {real, imag} */,
  {32'h44393126, 32'hc2af20d6} /* (14, 13, 30) {real, imag} */,
  {32'h42ecfbd2, 32'h4236ec18} /* (14, 13, 29) {real, imag} */,
  {32'hc2f5cd9f, 32'h43497a28} /* (14, 13, 28) {real, imag} */,
  {32'h42dca137, 32'hc31f0dc0} /* (14, 13, 27) {real, imag} */,
  {32'h42466eb3, 32'hc29e0a90} /* (14, 13, 26) {real, imag} */,
  {32'hc10f6bb8, 32'h4128ae5c} /* (14, 13, 25) {real, imag} */,
  {32'h428f7371, 32'h41e0f2dd} /* (14, 13, 24) {real, imag} */,
  {32'hc20f4eef, 32'h429d5259} /* (14, 13, 23) {real, imag} */,
  {32'h423c330f, 32'h40f6a368} /* (14, 13, 22) {real, imag} */,
  {32'h42501ad6, 32'hc31ebb0e} /* (14, 13, 21) {real, imag} */,
  {32'hc2651ea2, 32'hc2b359aa} /* (14, 13, 20) {real, imag} */,
  {32'h41b0012b, 32'hc1b048c2} /* (14, 13, 19) {real, imag} */,
  {32'hc21d72f4, 32'hc2a9aca4} /* (14, 13, 18) {real, imag} */,
  {32'hc13777b0, 32'h402ee158} /* (14, 13, 17) {real, imag} */,
  {32'h421cd716, 32'h00000000} /* (14, 13, 16) {real, imag} */,
  {32'hc13777b0, 32'hc02ee158} /* (14, 13, 15) {real, imag} */,
  {32'hc21d72f4, 32'h42a9aca4} /* (14, 13, 14) {real, imag} */,
  {32'h41b0012b, 32'h41b048c2} /* (14, 13, 13) {real, imag} */,
  {32'hc2651ea2, 32'h42b359aa} /* (14, 13, 12) {real, imag} */,
  {32'h42501ad6, 32'h431ebb0e} /* (14, 13, 11) {real, imag} */,
  {32'h423c330f, 32'hc0f6a368} /* (14, 13, 10) {real, imag} */,
  {32'hc20f4eef, 32'hc29d5259} /* (14, 13, 9) {real, imag} */,
  {32'h428f7371, 32'hc1e0f2dd} /* (14, 13, 8) {real, imag} */,
  {32'hc10f6bb8, 32'hc128ae5c} /* (14, 13, 7) {real, imag} */,
  {32'h42466eb3, 32'h429e0a90} /* (14, 13, 6) {real, imag} */,
  {32'h42dca137, 32'h431f0dc0} /* (14, 13, 5) {real, imag} */,
  {32'hc2f5cd9f, 32'hc3497a28} /* (14, 13, 4) {real, imag} */,
  {32'h42ecfbd2, 32'hc236ec18} /* (14, 13, 3) {real, imag} */,
  {32'h44393126, 32'h42af20d6} /* (14, 13, 2) {real, imag} */,
  {32'hc50c7100, 32'hc356be92} /* (14, 13, 1) {real, imag} */,
  {32'hc48fc6f2, 32'h00000000} /* (14, 13, 0) {real, imag} */,
  {32'hc4e09d72, 32'h435ab408} /* (14, 12, 31) {real, imag} */,
  {32'h441d5295, 32'hc08f8c40} /* (14, 12, 30) {real, imag} */,
  {32'h420fff30, 32'hc0a3fe78} /* (14, 12, 29) {real, imag} */,
  {32'hc3368df8, 32'h435ded6f} /* (14, 12, 28) {real, imag} */,
  {32'h436b0b42, 32'hc334201e} /* (14, 12, 27) {real, imag} */,
  {32'h423ff080, 32'hc07647a0} /* (14, 12, 26) {real, imag} */,
  {32'h42b62d54, 32'hc2827786} /* (14, 12, 25) {real, imag} */,
  {32'h429b0696, 32'hc12b286c} /* (14, 12, 24) {real, imag} */,
  {32'hc03fa6f0, 32'h41b25f66} /* (14, 12, 23) {real, imag} */,
  {32'h41300410, 32'hc24c06d3} /* (14, 12, 22) {real, imag} */,
  {32'h426293a6, 32'hc296cd13} /* (14, 12, 21) {real, imag} */,
  {32'hc19e270a, 32'hc2752baa} /* (14, 12, 20) {real, imag} */,
  {32'h423b815e, 32'h4206b4af} /* (14, 12, 19) {real, imag} */,
  {32'h41f64df0, 32'h4096a140} /* (14, 12, 18) {real, imag} */,
  {32'h41b43c5a, 32'hc2626c14} /* (14, 12, 17) {real, imag} */,
  {32'hc2b13818, 32'h00000000} /* (14, 12, 16) {real, imag} */,
  {32'h41b43c5a, 32'h42626c14} /* (14, 12, 15) {real, imag} */,
  {32'h41f64df0, 32'hc096a140} /* (14, 12, 14) {real, imag} */,
  {32'h423b815e, 32'hc206b4af} /* (14, 12, 13) {real, imag} */,
  {32'hc19e270a, 32'h42752baa} /* (14, 12, 12) {real, imag} */,
  {32'h426293a6, 32'h4296cd13} /* (14, 12, 11) {real, imag} */,
  {32'h41300410, 32'h424c06d3} /* (14, 12, 10) {real, imag} */,
  {32'hc03fa6f0, 32'hc1b25f66} /* (14, 12, 9) {real, imag} */,
  {32'h429b0696, 32'h412b286c} /* (14, 12, 8) {real, imag} */,
  {32'h42b62d54, 32'h42827786} /* (14, 12, 7) {real, imag} */,
  {32'h423ff080, 32'h407647a0} /* (14, 12, 6) {real, imag} */,
  {32'h436b0b42, 32'h4334201e} /* (14, 12, 5) {real, imag} */,
  {32'hc3368df8, 32'hc35ded6f} /* (14, 12, 4) {real, imag} */,
  {32'h420fff30, 32'h40a3fe78} /* (14, 12, 3) {real, imag} */,
  {32'h441d5295, 32'h408f8c40} /* (14, 12, 2) {real, imag} */,
  {32'hc4e09d72, 32'hc35ab408} /* (14, 12, 1) {real, imag} */,
  {32'hc414aa94, 32'h00000000} /* (14, 12, 0) {real, imag} */,
  {32'hc46d4421, 32'h42faf5f0} /* (14, 11, 31) {real, imag} */,
  {32'h440dd2ef, 32'h42a52262} /* (14, 11, 30) {real, imag} */,
  {32'h424b0bda, 32'h42626dce} /* (14, 11, 29) {real, imag} */,
  {32'hc2857418, 32'h42af0d4a} /* (14, 11, 28) {real, imag} */,
  {32'h42d2d22f, 32'hc31f544c} /* (14, 11, 27) {real, imag} */,
  {32'h429a83ac, 32'h41e74e43} /* (14, 11, 26) {real, imag} */,
  {32'hc28b99bd, 32'hc2dac313} /* (14, 11, 25) {real, imag} */,
  {32'h423fcbde, 32'hc1f83e0f} /* (14, 11, 24) {real, imag} */,
  {32'hc2edfb2e, 32'hc2d7caaf} /* (14, 11, 23) {real, imag} */,
  {32'hc2c22a4a, 32'hc235f358} /* (14, 11, 22) {real, imag} */,
  {32'hc29dc13e, 32'hc211af48} /* (14, 11, 21) {real, imag} */,
  {32'hc00b293c, 32'h4329155c} /* (14, 11, 20) {real, imag} */,
  {32'h42e1ed59, 32'h42223fa0} /* (14, 11, 19) {real, imag} */,
  {32'h427ad0ca, 32'h4131c800} /* (14, 11, 18) {real, imag} */,
  {32'h425e0d28, 32'h40397cc0} /* (14, 11, 17) {real, imag} */,
  {32'hc1b6b172, 32'h00000000} /* (14, 11, 16) {real, imag} */,
  {32'h425e0d28, 32'hc0397cc0} /* (14, 11, 15) {real, imag} */,
  {32'h427ad0ca, 32'hc131c800} /* (14, 11, 14) {real, imag} */,
  {32'h42e1ed59, 32'hc2223fa0} /* (14, 11, 13) {real, imag} */,
  {32'hc00b293c, 32'hc329155c} /* (14, 11, 12) {real, imag} */,
  {32'hc29dc13e, 32'h4211af48} /* (14, 11, 11) {real, imag} */,
  {32'hc2c22a4a, 32'h4235f358} /* (14, 11, 10) {real, imag} */,
  {32'hc2edfb2e, 32'h42d7caaf} /* (14, 11, 9) {real, imag} */,
  {32'h423fcbde, 32'h41f83e0f} /* (14, 11, 8) {real, imag} */,
  {32'hc28b99bd, 32'h42dac313} /* (14, 11, 7) {real, imag} */,
  {32'h429a83ac, 32'hc1e74e43} /* (14, 11, 6) {real, imag} */,
  {32'h42d2d22f, 32'h431f544c} /* (14, 11, 5) {real, imag} */,
  {32'hc2857418, 32'hc2af0d4a} /* (14, 11, 4) {real, imag} */,
  {32'h424b0bda, 32'hc2626dce} /* (14, 11, 3) {real, imag} */,
  {32'h440dd2ef, 32'hc2a52262} /* (14, 11, 2) {real, imag} */,
  {32'hc46d4421, 32'hc2faf5f0} /* (14, 11, 1) {real, imag} */,
  {32'h400f9e00, 32'h00000000} /* (14, 11, 0) {real, imag} */,
  {32'h4403599a, 32'hc37ad559} /* (14, 10, 31) {real, imag} */,
  {32'h428a6928, 32'h42ee1b4c} /* (14, 10, 30) {real, imag} */,
  {32'h421ef388, 32'h42665443} /* (14, 10, 29) {real, imag} */,
  {32'hc23a6c80, 32'hc0c2a070} /* (14, 10, 28) {real, imag} */,
  {32'hc347ac70, 32'h4273c50b} /* (14, 10, 27) {real, imag} */,
  {32'hc22420fc, 32'h42893e8c} /* (14, 10, 26) {real, imag} */,
  {32'hc2afe03b, 32'h41f93aed} /* (14, 10, 25) {real, imag} */,
  {32'h41cc75af, 32'h420df6d0} /* (14, 10, 24) {real, imag} */,
  {32'h411a8ba0, 32'h42f26aba} /* (14, 10, 23) {real, imag} */,
  {32'h41e793e2, 32'hc1343a3c} /* (14, 10, 22) {real, imag} */,
  {32'h40eaf9f0, 32'hc2901522} /* (14, 10, 21) {real, imag} */,
  {32'h426a1244, 32'hc201fbac} /* (14, 10, 20) {real, imag} */,
  {32'hc17845fa, 32'hc2fcaa9d} /* (14, 10, 19) {real, imag} */,
  {32'hc2f70479, 32'hc1d6fa10} /* (14, 10, 18) {real, imag} */,
  {32'hc2d7a252, 32'hc23f3dc0} /* (14, 10, 17) {real, imag} */,
  {32'hc18e3884, 32'h00000000} /* (14, 10, 16) {real, imag} */,
  {32'hc2d7a252, 32'h423f3dc0} /* (14, 10, 15) {real, imag} */,
  {32'hc2f70479, 32'h41d6fa10} /* (14, 10, 14) {real, imag} */,
  {32'hc17845fa, 32'h42fcaa9d} /* (14, 10, 13) {real, imag} */,
  {32'h426a1244, 32'h4201fbac} /* (14, 10, 12) {real, imag} */,
  {32'h40eaf9f0, 32'h42901522} /* (14, 10, 11) {real, imag} */,
  {32'h41e793e2, 32'h41343a3c} /* (14, 10, 10) {real, imag} */,
  {32'h411a8ba0, 32'hc2f26aba} /* (14, 10, 9) {real, imag} */,
  {32'h41cc75af, 32'hc20df6d0} /* (14, 10, 8) {real, imag} */,
  {32'hc2afe03b, 32'hc1f93aed} /* (14, 10, 7) {real, imag} */,
  {32'hc22420fc, 32'hc2893e8c} /* (14, 10, 6) {real, imag} */,
  {32'hc347ac70, 32'hc273c50b} /* (14, 10, 5) {real, imag} */,
  {32'hc23a6c80, 32'h40c2a070} /* (14, 10, 4) {real, imag} */,
  {32'h421ef388, 32'hc2665443} /* (14, 10, 3) {real, imag} */,
  {32'h428a6928, 32'hc2ee1b4c} /* (14, 10, 2) {real, imag} */,
  {32'h4403599a, 32'h437ad559} /* (14, 10, 1) {real, imag} */,
  {32'h447a318d, 32'h00000000} /* (14, 10, 0) {real, imag} */,
  {32'h449e886a, 32'hc3e28374} /* (14, 9, 31) {real, imag} */,
  {32'hc3f0dde2, 32'h4349d9ac} /* (14, 9, 30) {real, imag} */,
  {32'hc1afbbfa, 32'h4321b840} /* (14, 9, 29) {real, imag} */,
  {32'hc20afe17, 32'hc07f2720} /* (14, 9, 28) {real, imag} */,
  {32'hc3372b78, 32'h4371d200} /* (14, 9, 27) {real, imag} */,
  {32'h428a7a96, 32'hc1bdea17} /* (14, 9, 26) {real, imag} */,
  {32'hc2ea040f, 32'hc0ebb558} /* (14, 9, 25) {real, imag} */,
  {32'h419a98d6, 32'h42e55cfa} /* (14, 9, 24) {real, imag} */,
  {32'hbfb7df40, 32'h41becc8a} /* (14, 9, 23) {real, imag} */,
  {32'h419865b4, 32'h4293d302} /* (14, 9, 22) {real, imag} */,
  {32'hc19b3667, 32'h42ae5b31} /* (14, 9, 21) {real, imag} */,
  {32'h42efff5a, 32'hc24f89c3} /* (14, 9, 20) {real, imag} */,
  {32'hc1d3a997, 32'hc2886278} /* (14, 9, 19) {real, imag} */,
  {32'hc1d4cf1e, 32'h42b0bfff} /* (14, 9, 18) {real, imag} */,
  {32'h428ca143, 32'hc257fc94} /* (14, 9, 17) {real, imag} */,
  {32'h41eb7177, 32'h00000000} /* (14, 9, 16) {real, imag} */,
  {32'h428ca143, 32'h4257fc94} /* (14, 9, 15) {real, imag} */,
  {32'hc1d4cf1e, 32'hc2b0bfff} /* (14, 9, 14) {real, imag} */,
  {32'hc1d3a997, 32'h42886278} /* (14, 9, 13) {real, imag} */,
  {32'h42efff5a, 32'h424f89c3} /* (14, 9, 12) {real, imag} */,
  {32'hc19b3667, 32'hc2ae5b31} /* (14, 9, 11) {real, imag} */,
  {32'h419865b4, 32'hc293d302} /* (14, 9, 10) {real, imag} */,
  {32'hbfb7df40, 32'hc1becc8a} /* (14, 9, 9) {real, imag} */,
  {32'h419a98d6, 32'hc2e55cfa} /* (14, 9, 8) {real, imag} */,
  {32'hc2ea040f, 32'h40ebb558} /* (14, 9, 7) {real, imag} */,
  {32'h428a7a96, 32'h41bdea17} /* (14, 9, 6) {real, imag} */,
  {32'hc3372b78, 32'hc371d200} /* (14, 9, 5) {real, imag} */,
  {32'hc20afe17, 32'h407f2720} /* (14, 9, 4) {real, imag} */,
  {32'hc1afbbfa, 32'hc321b840} /* (14, 9, 3) {real, imag} */,
  {32'hc3f0dde2, 32'hc349d9ac} /* (14, 9, 2) {real, imag} */,
  {32'h449e886a, 32'h43e28374} /* (14, 9, 1) {real, imag} */,
  {32'h44db576a, 32'h00000000} /* (14, 9, 0) {real, imag} */,
  {32'h44c06eed, 32'hc408687f} /* (14, 8, 31) {real, imag} */,
  {32'hc42836ce, 32'h43c824d8} /* (14, 8, 30) {real, imag} */,
  {32'hc232e6fd, 32'h42fede0a} /* (14, 8, 29) {real, imag} */,
  {32'h430faa86, 32'hc27f856b} /* (14, 8, 28) {real, imag} */,
  {32'hc2abe6b2, 32'h40b39e60} /* (14, 8, 27) {real, imag} */,
  {32'h415966e8, 32'h42e50d74} /* (14, 8, 26) {real, imag} */,
  {32'hc25734cc, 32'h42c0bca1} /* (14, 8, 25) {real, imag} */,
  {32'hc2af2586, 32'h42d209e0} /* (14, 8, 24) {real, imag} */,
  {32'hc28abefe, 32'hc26f2a16} /* (14, 8, 23) {real, imag} */,
  {32'hc24d49ce, 32'hc2b2ff1a} /* (14, 8, 22) {real, imag} */,
  {32'hc24a0bce, 32'hc1cf3890} /* (14, 8, 21) {real, imag} */,
  {32'hc24dcb82, 32'h41995ce4} /* (14, 8, 20) {real, imag} */,
  {32'h428d5b78, 32'hc1d6a109} /* (14, 8, 19) {real, imag} */,
  {32'hc2662a72, 32'h429bf8b8} /* (14, 8, 18) {real, imag} */,
  {32'hc2ae477e, 32'h42d6a18a} /* (14, 8, 17) {real, imag} */,
  {32'h40dac844, 32'h00000000} /* (14, 8, 16) {real, imag} */,
  {32'hc2ae477e, 32'hc2d6a18a} /* (14, 8, 15) {real, imag} */,
  {32'hc2662a72, 32'hc29bf8b8} /* (14, 8, 14) {real, imag} */,
  {32'h428d5b78, 32'h41d6a109} /* (14, 8, 13) {real, imag} */,
  {32'hc24dcb82, 32'hc1995ce4} /* (14, 8, 12) {real, imag} */,
  {32'hc24a0bce, 32'h41cf3890} /* (14, 8, 11) {real, imag} */,
  {32'hc24d49ce, 32'h42b2ff1a} /* (14, 8, 10) {real, imag} */,
  {32'hc28abefe, 32'h426f2a16} /* (14, 8, 9) {real, imag} */,
  {32'hc2af2586, 32'hc2d209e0} /* (14, 8, 8) {real, imag} */,
  {32'hc25734cc, 32'hc2c0bca1} /* (14, 8, 7) {real, imag} */,
  {32'h415966e8, 32'hc2e50d74} /* (14, 8, 6) {real, imag} */,
  {32'hc2abe6b2, 32'hc0b39e60} /* (14, 8, 5) {real, imag} */,
  {32'h430faa86, 32'h427f856b} /* (14, 8, 4) {real, imag} */,
  {32'hc232e6fd, 32'hc2fede0a} /* (14, 8, 3) {real, imag} */,
  {32'hc42836ce, 32'hc3c824d8} /* (14, 8, 2) {real, imag} */,
  {32'h44c06eed, 32'h4408687f} /* (14, 8, 1) {real, imag} */,
  {32'h45025d86, 32'h00000000} /* (14, 8, 0) {real, imag} */,
  {32'h44dac22e, 32'hc42ce0dc} /* (14, 7, 31) {real, imag} */,
  {32'hc43d8a21, 32'h43d09a10} /* (14, 7, 30) {real, imag} */,
  {32'hc27d79b9, 32'h427bc146} /* (14, 7, 29) {real, imag} */,
  {32'h431e7320, 32'hc2a33d59} /* (14, 7, 28) {real, imag} */,
  {32'hc2f87f3b, 32'h41c52d24} /* (14, 7, 27) {real, imag} */,
  {32'h424ca9ca, 32'h42c65d18} /* (14, 7, 26) {real, imag} */,
  {32'hc2308158, 32'h41160ef8} /* (14, 7, 25) {real, imag} */,
  {32'hc2ef662a, 32'hc1e13010} /* (14, 7, 24) {real, imag} */,
  {32'hc1c20a0c, 32'h4284587a} /* (14, 7, 23) {real, imag} */,
  {32'h4233457d, 32'hc2d10b04} /* (14, 7, 22) {real, imag} */,
  {32'hc29feb72, 32'h41ba1fb4} /* (14, 7, 21) {real, imag} */,
  {32'h41ec90a1, 32'hc21e08d2} /* (14, 7, 20) {real, imag} */,
  {32'h42432c82, 32'hc292cdee} /* (14, 7, 19) {real, imag} */,
  {32'hc19034ce, 32'h42a9f644} /* (14, 7, 18) {real, imag} */,
  {32'h41185129, 32'h421ec9e6} /* (14, 7, 17) {real, imag} */,
  {32'h42c48baa, 32'h00000000} /* (14, 7, 16) {real, imag} */,
  {32'h41185129, 32'hc21ec9e6} /* (14, 7, 15) {real, imag} */,
  {32'hc19034ce, 32'hc2a9f644} /* (14, 7, 14) {real, imag} */,
  {32'h42432c82, 32'h4292cdee} /* (14, 7, 13) {real, imag} */,
  {32'h41ec90a1, 32'h421e08d2} /* (14, 7, 12) {real, imag} */,
  {32'hc29feb72, 32'hc1ba1fb4} /* (14, 7, 11) {real, imag} */,
  {32'h4233457d, 32'h42d10b04} /* (14, 7, 10) {real, imag} */,
  {32'hc1c20a0c, 32'hc284587a} /* (14, 7, 9) {real, imag} */,
  {32'hc2ef662a, 32'h41e13010} /* (14, 7, 8) {real, imag} */,
  {32'hc2308158, 32'hc1160ef8} /* (14, 7, 7) {real, imag} */,
  {32'h424ca9ca, 32'hc2c65d18} /* (14, 7, 6) {real, imag} */,
  {32'hc2f87f3b, 32'hc1c52d24} /* (14, 7, 5) {real, imag} */,
  {32'h431e7320, 32'h42a33d59} /* (14, 7, 4) {real, imag} */,
  {32'hc27d79b9, 32'hc27bc146} /* (14, 7, 3) {real, imag} */,
  {32'hc43d8a21, 32'hc3d09a10} /* (14, 7, 2) {real, imag} */,
  {32'h44dac22e, 32'h442ce0dc} /* (14, 7, 1) {real, imag} */,
  {32'h451048ba, 32'h00000000} /* (14, 7, 0) {real, imag} */,
  {32'h44eda8a1, 32'hc47e9606} /* (14, 6, 31) {real, imag} */,
  {32'hc4211a33, 32'h440561f6} /* (14, 6, 30) {real, imag} */,
  {32'hc2e5971d, 32'h42dfb66a} /* (14, 6, 29) {real, imag} */,
  {32'h42df21a4, 32'h40f10030} /* (14, 6, 28) {real, imag} */,
  {32'hc3298158, 32'h432bdf27} /* (14, 6, 27) {real, imag} */,
  {32'h42b020ac, 32'h41460510} /* (14, 6, 26) {real, imag} */,
  {32'h424da6f0, 32'hc309a9f4} /* (14, 6, 25) {real, imag} */,
  {32'h417e1684, 32'h41398c02} /* (14, 6, 24) {real, imag} */,
  {32'hbfa09f80, 32'h42da7bcd} /* (14, 6, 23) {real, imag} */,
  {32'h429e5e76, 32'h42543b9c} /* (14, 6, 22) {real, imag} */,
  {32'hc1b83994, 32'h42e6096f} /* (14, 6, 21) {real, imag} */,
  {32'h41b1b446, 32'h425f9f6c} /* (14, 6, 20) {real, imag} */,
  {32'hc2b2b89d, 32'h416b60be} /* (14, 6, 19) {real, imag} */,
  {32'hc24181c4, 32'hc2161255} /* (14, 6, 18) {real, imag} */,
  {32'hc252aace, 32'hc29db1f6} /* (14, 6, 17) {real, imag} */,
  {32'hc28a7e99, 32'h00000000} /* (14, 6, 16) {real, imag} */,
  {32'hc252aace, 32'h429db1f6} /* (14, 6, 15) {real, imag} */,
  {32'hc24181c4, 32'h42161255} /* (14, 6, 14) {real, imag} */,
  {32'hc2b2b89d, 32'hc16b60be} /* (14, 6, 13) {real, imag} */,
  {32'h41b1b446, 32'hc25f9f6c} /* (14, 6, 12) {real, imag} */,
  {32'hc1b83994, 32'hc2e6096f} /* (14, 6, 11) {real, imag} */,
  {32'h429e5e76, 32'hc2543b9c} /* (14, 6, 10) {real, imag} */,
  {32'hbfa09f80, 32'hc2da7bcd} /* (14, 6, 9) {real, imag} */,
  {32'h417e1684, 32'hc1398c02} /* (14, 6, 8) {real, imag} */,
  {32'h424da6f0, 32'h4309a9f4} /* (14, 6, 7) {real, imag} */,
  {32'h42b020ac, 32'hc1460510} /* (14, 6, 6) {real, imag} */,
  {32'hc3298158, 32'hc32bdf27} /* (14, 6, 5) {real, imag} */,
  {32'h42df21a4, 32'hc0f10030} /* (14, 6, 4) {real, imag} */,
  {32'hc2e5971d, 32'hc2dfb66a} /* (14, 6, 3) {real, imag} */,
  {32'hc4211a33, 32'hc40561f6} /* (14, 6, 2) {real, imag} */,
  {32'h44eda8a1, 32'h447e9606} /* (14, 6, 1) {real, imag} */,
  {32'h451cdc75, 32'h00000000} /* (14, 6, 0) {real, imag} */,
  {32'h44dfb27e, 32'hc4d1b090} /* (14, 5, 31) {real, imag} */,
  {32'hc3479b68, 32'h4428d9a4} /* (14, 5, 30) {real, imag} */,
  {32'hc2b9cbd8, 32'h4311dee0} /* (14, 5, 29) {real, imag} */,
  {32'hc31009a2, 32'hc101b930} /* (14, 5, 28) {real, imag} */,
  {32'hc3428f38, 32'h421708a6} /* (14, 5, 27) {real, imag} */,
  {32'h42c2df88, 32'h42e4e47c} /* (14, 5, 26) {real, imag} */,
  {32'hc2c38458, 32'hc25046ca} /* (14, 5, 25) {real, imag} */,
  {32'h426b4070, 32'hc152bf00} /* (14, 5, 24) {real, imag} */,
  {32'hc2705a16, 32'hc2186c1c} /* (14, 5, 23) {real, imag} */,
  {32'hc0c94938, 32'hc27b4933} /* (14, 5, 22) {real, imag} */,
  {32'hc1ae2e09, 32'h420d2f50} /* (14, 5, 21) {real, imag} */,
  {32'h42969e64, 32'h4047c7e8} /* (14, 5, 20) {real, imag} */,
  {32'h41ccb077, 32'h40f2613c} /* (14, 5, 19) {real, imag} */,
  {32'hc172ceb8, 32'h419e443c} /* (14, 5, 18) {real, imag} */,
  {32'h414d447c, 32'h428c892f} /* (14, 5, 17) {real, imag} */,
  {32'h422b1444, 32'h00000000} /* (14, 5, 16) {real, imag} */,
  {32'h414d447c, 32'hc28c892f} /* (14, 5, 15) {real, imag} */,
  {32'hc172ceb8, 32'hc19e443c} /* (14, 5, 14) {real, imag} */,
  {32'h41ccb077, 32'hc0f2613c} /* (14, 5, 13) {real, imag} */,
  {32'h42969e64, 32'hc047c7e8} /* (14, 5, 12) {real, imag} */,
  {32'hc1ae2e09, 32'hc20d2f50} /* (14, 5, 11) {real, imag} */,
  {32'hc0c94938, 32'h427b4933} /* (14, 5, 10) {real, imag} */,
  {32'hc2705a16, 32'h42186c1c} /* (14, 5, 9) {real, imag} */,
  {32'h426b4070, 32'h4152bf00} /* (14, 5, 8) {real, imag} */,
  {32'hc2c38458, 32'h425046ca} /* (14, 5, 7) {real, imag} */,
  {32'h42c2df88, 32'hc2e4e47c} /* (14, 5, 6) {real, imag} */,
  {32'hc3428f38, 32'hc21708a6} /* (14, 5, 5) {real, imag} */,
  {32'hc31009a2, 32'h4101b930} /* (14, 5, 4) {real, imag} */,
  {32'hc2b9cbd8, 32'hc311dee0} /* (14, 5, 3) {real, imag} */,
  {32'hc3479b68, 32'hc428d9a4} /* (14, 5, 2) {real, imag} */,
  {32'h44dfb27e, 32'h44d1b090} /* (14, 5, 1) {real, imag} */,
  {32'h451d2969, 32'h00000000} /* (14, 5, 0) {real, imag} */,
  {32'h44c8f5de, 32'hc5040571} /* (14, 4, 31) {real, imag} */,
  {32'h426d3e18, 32'h44377415} /* (14, 4, 30) {real, imag} */,
  {32'hc2a543b5, 32'h4343dbb2} /* (14, 4, 29) {real, imag} */,
  {32'hc3534e22, 32'h3fb23b20} /* (14, 4, 28) {real, imag} */,
  {32'hc3459586, 32'h41c9647c} /* (14, 4, 27) {real, imag} */,
  {32'h42b73499, 32'h42b96754} /* (14, 4, 26) {real, imag} */,
  {32'hc31c706b, 32'hc1a69350} /* (14, 4, 25) {real, imag} */,
  {32'h41345489, 32'hc1836e42} /* (14, 4, 24) {real, imag} */,
  {32'h40f40c78, 32'hc18d2958} /* (14, 4, 23) {real, imag} */,
  {32'hc224fc52, 32'h418c299a} /* (14, 4, 22) {real, imag} */,
  {32'hc2143a9c, 32'hc1e5cd5b} /* (14, 4, 21) {real, imag} */,
  {32'h41c36ac2, 32'hc174fe4a} /* (14, 4, 20) {real, imag} */,
  {32'h4214524a, 32'h41077ee0} /* (14, 4, 19) {real, imag} */,
  {32'hc1ab4774, 32'h419f87c0} /* (14, 4, 18) {real, imag} */,
  {32'h40815148, 32'hc14b6e30} /* (14, 4, 17) {real, imag} */,
  {32'h428163af, 32'h00000000} /* (14, 4, 16) {real, imag} */,
  {32'h40815148, 32'h414b6e30} /* (14, 4, 15) {real, imag} */,
  {32'hc1ab4774, 32'hc19f87c0} /* (14, 4, 14) {real, imag} */,
  {32'h4214524a, 32'hc1077ee0} /* (14, 4, 13) {real, imag} */,
  {32'h41c36ac2, 32'h4174fe4a} /* (14, 4, 12) {real, imag} */,
  {32'hc2143a9c, 32'h41e5cd5b} /* (14, 4, 11) {real, imag} */,
  {32'hc224fc52, 32'hc18c299a} /* (14, 4, 10) {real, imag} */,
  {32'h40f40c78, 32'h418d2958} /* (14, 4, 9) {real, imag} */,
  {32'h41345489, 32'h41836e42} /* (14, 4, 8) {real, imag} */,
  {32'hc31c706b, 32'h41a69350} /* (14, 4, 7) {real, imag} */,
  {32'h42b73499, 32'hc2b96754} /* (14, 4, 6) {real, imag} */,
  {32'hc3459586, 32'hc1c9647c} /* (14, 4, 5) {real, imag} */,
  {32'hc3534e22, 32'hbfb23b20} /* (14, 4, 4) {real, imag} */,
  {32'hc2a543b5, 32'hc343dbb2} /* (14, 4, 3) {real, imag} */,
  {32'h426d3e18, 32'hc4377415} /* (14, 4, 2) {real, imag} */,
  {32'h44c8f5de, 32'h45040571} /* (14, 4, 1) {real, imag} */,
  {32'h45355c83, 32'h00000000} /* (14, 4, 0) {real, imag} */,
  {32'h44c4a16e, 32'hc507d3bd} /* (14, 3, 31) {real, imag} */,
  {32'h42b1c7c0, 32'h443fc5b2} /* (14, 3, 30) {real, imag} */,
  {32'hc3270b19, 32'h428da4a8} /* (14, 3, 29) {real, imag} */,
  {32'hc3049aba, 32'h42a92cb4} /* (14, 3, 28) {real, imag} */,
  {32'hc2fc6796, 32'hc28562de} /* (14, 3, 27) {real, imag} */,
  {32'h42b61db6, 32'hc1375401} /* (14, 3, 26) {real, imag} */,
  {32'h42b03496, 32'hc301f9f0} /* (14, 3, 25) {real, imag} */,
  {32'h4168fd13, 32'hc247012a} /* (14, 3, 24) {real, imag} */,
  {32'hc131e2c8, 32'hc2740987} /* (14, 3, 23) {real, imag} */,
  {32'hc29caf82, 32'hc1bed3de} /* (14, 3, 22) {real, imag} */,
  {32'hc22b96ea, 32'h423c0677} /* (14, 3, 21) {real, imag} */,
  {32'h40b7bbc0, 32'hc1ec4857} /* (14, 3, 20) {real, imag} */,
  {32'h41af3d94, 32'hc1654424} /* (14, 3, 19) {real, imag} */,
  {32'h426fc812, 32'hc2b02cad} /* (14, 3, 18) {real, imag} */,
  {32'hc3071082, 32'h4265ebd8} /* (14, 3, 17) {real, imag} */,
  {32'h410658bc, 32'h00000000} /* (14, 3, 16) {real, imag} */,
  {32'hc3071082, 32'hc265ebd8} /* (14, 3, 15) {real, imag} */,
  {32'h426fc812, 32'h42b02cad} /* (14, 3, 14) {real, imag} */,
  {32'h41af3d94, 32'h41654424} /* (14, 3, 13) {real, imag} */,
  {32'h40b7bbc0, 32'h41ec4857} /* (14, 3, 12) {real, imag} */,
  {32'hc22b96ea, 32'hc23c0677} /* (14, 3, 11) {real, imag} */,
  {32'hc29caf82, 32'h41bed3de} /* (14, 3, 10) {real, imag} */,
  {32'hc131e2c8, 32'h42740987} /* (14, 3, 9) {real, imag} */,
  {32'h4168fd13, 32'h4247012a} /* (14, 3, 8) {real, imag} */,
  {32'h42b03496, 32'h4301f9f0} /* (14, 3, 7) {real, imag} */,
  {32'h42b61db6, 32'h41375401} /* (14, 3, 6) {real, imag} */,
  {32'hc2fc6796, 32'h428562de} /* (14, 3, 5) {real, imag} */,
  {32'hc3049aba, 32'hc2a92cb4} /* (14, 3, 4) {real, imag} */,
  {32'hc3270b19, 32'hc28da4a8} /* (14, 3, 3) {real, imag} */,
  {32'h42b1c7c0, 32'hc43fc5b2} /* (14, 3, 2) {real, imag} */,
  {32'h44c4a16e, 32'h4507d3bd} /* (14, 3, 1) {real, imag} */,
  {32'h4541208e, 32'h00000000} /* (14, 3, 0) {real, imag} */,
  {32'h44c9cfd6, 32'hc5020043} /* (14, 2, 31) {real, imag} */,
  {32'h4332b0cc, 32'h4429c3ce} /* (14, 2, 30) {real, imag} */,
  {32'hc2af7afe, 32'h42f53f8e} /* (14, 2, 29) {real, imag} */,
  {32'hc2af48ee, 32'h4316ea52} /* (14, 2, 28) {real, imag} */,
  {32'hc368f1f9, 32'hc28f14d2} /* (14, 2, 27) {real, imag} */,
  {32'hc28879c2, 32'hc2055982} /* (14, 2, 26) {real, imag} */,
  {32'hc24d95b9, 32'hc2f4e82c} /* (14, 2, 25) {real, imag} */,
  {32'hc2017459, 32'hc29e04d4} /* (14, 2, 24) {real, imag} */,
  {32'h41fffc18, 32'hc2f63932} /* (14, 2, 23) {real, imag} */,
  {32'hc2824dd6, 32'h42921c43} /* (14, 2, 22) {real, imag} */,
  {32'hc26f0c84, 32'hc21945ca} /* (14, 2, 21) {real, imag} */,
  {32'h426ebd4e, 32'h4270a07f} /* (14, 2, 20) {real, imag} */,
  {32'hc28a6c88, 32'h42154fa8} /* (14, 2, 19) {real, imag} */,
  {32'h41571d22, 32'h42c832b4} /* (14, 2, 18) {real, imag} */,
  {32'hc14fa020, 32'hc210795c} /* (14, 2, 17) {real, imag} */,
  {32'h4200a05f, 32'h00000000} /* (14, 2, 16) {real, imag} */,
  {32'hc14fa020, 32'h4210795c} /* (14, 2, 15) {real, imag} */,
  {32'h41571d22, 32'hc2c832b4} /* (14, 2, 14) {real, imag} */,
  {32'hc28a6c88, 32'hc2154fa8} /* (14, 2, 13) {real, imag} */,
  {32'h426ebd4e, 32'hc270a07f} /* (14, 2, 12) {real, imag} */,
  {32'hc26f0c84, 32'h421945ca} /* (14, 2, 11) {real, imag} */,
  {32'hc2824dd6, 32'hc2921c43} /* (14, 2, 10) {real, imag} */,
  {32'h41fffc18, 32'h42f63932} /* (14, 2, 9) {real, imag} */,
  {32'hc2017459, 32'h429e04d4} /* (14, 2, 8) {real, imag} */,
  {32'hc24d95b9, 32'h42f4e82c} /* (14, 2, 7) {real, imag} */,
  {32'hc28879c2, 32'h42055982} /* (14, 2, 6) {real, imag} */,
  {32'hc368f1f9, 32'h428f14d2} /* (14, 2, 5) {real, imag} */,
  {32'hc2af48ee, 32'hc316ea52} /* (14, 2, 4) {real, imag} */,
  {32'hc2af7afe, 32'hc2f53f8e} /* (14, 2, 3) {real, imag} */,
  {32'h4332b0cc, 32'hc429c3ce} /* (14, 2, 2) {real, imag} */,
  {32'h44c9cfd6, 32'h45020043} /* (14, 2, 1) {real, imag} */,
  {32'h4532c1de, 32'h00000000} /* (14, 2, 0) {real, imag} */,
  {32'h44ce41bc, 32'hc5018ebb} /* (14, 1, 31) {real, imag} */,
  {32'h42d31b54, 32'h44098264} /* (14, 1, 30) {real, imag} */,
  {32'hc34dd37e, 32'h42adc47e} /* (14, 1, 29) {real, imag} */,
  {32'hc30b5042, 32'h42c5e3a7} /* (14, 1, 28) {real, imag} */,
  {32'hc31eb710, 32'hc289b560} /* (14, 1, 27) {real, imag} */,
  {32'hc229b154, 32'h4136a75c} /* (14, 1, 26) {real, imag} */,
  {32'hc2aa6b25, 32'h4263d979} /* (14, 1, 25) {real, imag} */,
  {32'h419c20bc, 32'h40894a34} /* (14, 1, 24) {real, imag} */,
  {32'h414e8518, 32'h40da920c} /* (14, 1, 23) {real, imag} */,
  {32'hc2984894, 32'hc2a82c32} /* (14, 1, 22) {real, imag} */,
  {32'hc251808e, 32'hc1619c5f} /* (14, 1, 21) {real, imag} */,
  {32'h424a32e9, 32'h4273bb48} /* (14, 1, 20) {real, imag} */,
  {32'h4208b679, 32'hc2c4ae75} /* (14, 1, 19) {real, imag} */,
  {32'h414f8b78, 32'h41c64800} /* (14, 1, 18) {real, imag} */,
  {32'h41e0dd57, 32'h42928cb8} /* (14, 1, 17) {real, imag} */,
  {32'h42047007, 32'h00000000} /* (14, 1, 16) {real, imag} */,
  {32'h41e0dd57, 32'hc2928cb8} /* (14, 1, 15) {real, imag} */,
  {32'h414f8b78, 32'hc1c64800} /* (14, 1, 14) {real, imag} */,
  {32'h4208b679, 32'h42c4ae75} /* (14, 1, 13) {real, imag} */,
  {32'h424a32e9, 32'hc273bb48} /* (14, 1, 12) {real, imag} */,
  {32'hc251808e, 32'h41619c5f} /* (14, 1, 11) {real, imag} */,
  {32'hc2984894, 32'h42a82c32} /* (14, 1, 10) {real, imag} */,
  {32'h414e8518, 32'hc0da920c} /* (14, 1, 9) {real, imag} */,
  {32'h419c20bc, 32'hc0894a34} /* (14, 1, 8) {real, imag} */,
  {32'hc2aa6b25, 32'hc263d979} /* (14, 1, 7) {real, imag} */,
  {32'hc229b154, 32'hc136a75c} /* (14, 1, 6) {real, imag} */,
  {32'hc31eb710, 32'h4289b560} /* (14, 1, 5) {real, imag} */,
  {32'hc30b5042, 32'hc2c5e3a7} /* (14, 1, 4) {real, imag} */,
  {32'hc34dd37e, 32'hc2adc47e} /* (14, 1, 3) {real, imag} */,
  {32'h42d31b54, 32'hc4098264} /* (14, 1, 2) {real, imag} */,
  {32'h44ce41bc, 32'h45018ebb} /* (14, 1, 1) {real, imag} */,
  {32'h4522cb82, 32'h00000000} /* (14, 1, 0) {real, imag} */,
  {32'h44d3fa4d, 32'hc4d42970} /* (14, 0, 31) {real, imag} */,
  {32'hc3073970, 32'h43be42ef} /* (14, 0, 30) {real, imag} */,
  {32'hc3097bba, 32'h41162d70} /* (14, 0, 29) {real, imag} */,
  {32'hc2e7c704, 32'h43077f51} /* (14, 0, 28) {real, imag} */,
  {32'hc2ffa789, 32'hc2326b57} /* (14, 0, 27) {real, imag} */,
  {32'h42300d59, 32'hc1953d26} /* (14, 0, 26) {real, imag} */,
  {32'h41da6579, 32'hc11552f1} /* (14, 0, 25) {real, imag} */,
  {32'hc133bee6, 32'hc2245811} /* (14, 0, 24) {real, imag} */,
  {32'hc260688e, 32'h4102426c} /* (14, 0, 23) {real, imag} */,
  {32'h414bb42c, 32'hc1fa18d4} /* (14, 0, 22) {real, imag} */,
  {32'h422b6e2d, 32'h424acfc9} /* (14, 0, 21) {real, imag} */,
  {32'hc0d3f4c6, 32'h4122cb10} /* (14, 0, 20) {real, imag} */,
  {32'h408b3bf8, 32'h41f94e1c} /* (14, 0, 19) {real, imag} */,
  {32'h4252c632, 32'hc2591080} /* (14, 0, 18) {real, imag} */,
  {32'hc230546c, 32'h4164105c} /* (14, 0, 17) {real, imag} */,
  {32'hc20b1247, 32'h00000000} /* (14, 0, 16) {real, imag} */,
  {32'hc230546c, 32'hc164105c} /* (14, 0, 15) {real, imag} */,
  {32'h4252c632, 32'h42591080} /* (14, 0, 14) {real, imag} */,
  {32'h408b3bf8, 32'hc1f94e1c} /* (14, 0, 13) {real, imag} */,
  {32'hc0d3f4c6, 32'hc122cb10} /* (14, 0, 12) {real, imag} */,
  {32'h422b6e2d, 32'hc24acfc9} /* (14, 0, 11) {real, imag} */,
  {32'h414bb42c, 32'h41fa18d4} /* (14, 0, 10) {real, imag} */,
  {32'hc260688e, 32'hc102426c} /* (14, 0, 9) {real, imag} */,
  {32'hc133bee6, 32'h42245811} /* (14, 0, 8) {real, imag} */,
  {32'h41da6579, 32'h411552f1} /* (14, 0, 7) {real, imag} */,
  {32'h42300d59, 32'h41953d26} /* (14, 0, 6) {real, imag} */,
  {32'hc2ffa789, 32'h42326b57} /* (14, 0, 5) {real, imag} */,
  {32'hc2e7c704, 32'hc3077f51} /* (14, 0, 4) {real, imag} */,
  {32'hc3097bba, 32'hc1162d70} /* (14, 0, 3) {real, imag} */,
  {32'hc3073970, 32'hc3be42ef} /* (14, 0, 2) {real, imag} */,
  {32'h44d3fa4d, 32'h44d42970} /* (14, 0, 1) {real, imag} */,
  {32'h45126baa, 32'h00000000} /* (14, 0, 0) {real, imag} */,
  {32'h453a3993, 32'hc4dc5cca} /* (13, 31, 31) {real, imag} */,
  {32'hc42e461c, 32'h43b3c684} /* (13, 31, 30) {real, imag} */,
  {32'hc2c73438, 32'h41a9777c} /* (13, 31, 29) {real, imag} */,
  {32'hc1e864d4, 32'hc1ad0c28} /* (13, 31, 28) {real, imag} */,
  {32'hc2e31f01, 32'hc30bf3d8} /* (13, 31, 27) {real, imag} */,
  {32'h4284e654, 32'hc2cdb984} /* (13, 31, 26) {real, imag} */,
  {32'hc1b513b2, 32'h423a7baa} /* (13, 31, 25) {real, imag} */,
  {32'hc29db974, 32'h41f60137} /* (13, 31, 24) {real, imag} */,
  {32'hc2c3b318, 32'h42bdd816} /* (13, 31, 23) {real, imag} */,
  {32'h3f4e1e20, 32'h4237fc3c} /* (13, 31, 22) {real, imag} */,
  {32'h40d13d94, 32'h423d02ab} /* (13, 31, 21) {real, imag} */,
  {32'hc09ed370, 32'hc18dddf2} /* (13, 31, 20) {real, imag} */,
  {32'hc20ca99c, 32'hc1af6db4} /* (13, 31, 19) {real, imag} */,
  {32'h421516be, 32'h426e6ce6} /* (13, 31, 18) {real, imag} */,
  {32'h41a8c7a0, 32'h4218a27e} /* (13, 31, 17) {real, imag} */,
  {32'h42392964, 32'h00000000} /* (13, 31, 16) {real, imag} */,
  {32'h41a8c7a0, 32'hc218a27e} /* (13, 31, 15) {real, imag} */,
  {32'h421516be, 32'hc26e6ce6} /* (13, 31, 14) {real, imag} */,
  {32'hc20ca99c, 32'h41af6db4} /* (13, 31, 13) {real, imag} */,
  {32'hc09ed370, 32'h418dddf2} /* (13, 31, 12) {real, imag} */,
  {32'h40d13d94, 32'hc23d02ab} /* (13, 31, 11) {real, imag} */,
  {32'h3f4e1e20, 32'hc237fc3c} /* (13, 31, 10) {real, imag} */,
  {32'hc2c3b318, 32'hc2bdd816} /* (13, 31, 9) {real, imag} */,
  {32'hc29db974, 32'hc1f60137} /* (13, 31, 8) {real, imag} */,
  {32'hc1b513b2, 32'hc23a7baa} /* (13, 31, 7) {real, imag} */,
  {32'h4284e654, 32'h42cdb984} /* (13, 31, 6) {real, imag} */,
  {32'hc2e31f01, 32'h430bf3d8} /* (13, 31, 5) {real, imag} */,
  {32'hc1e864d4, 32'h41ad0c28} /* (13, 31, 4) {real, imag} */,
  {32'hc2c73438, 32'hc1a9777c} /* (13, 31, 3) {real, imag} */,
  {32'hc42e461c, 32'hc3b3c684} /* (13, 31, 2) {real, imag} */,
  {32'h453a3993, 32'h44dc5cca} /* (13, 31, 1) {real, imag} */,
  {32'h45708aa0, 32'h00000000} /* (13, 31, 0) {real, imag} */,
  {32'h4554571a, 32'hc4abdc7e} /* (13, 30, 31) {real, imag} */,
  {32'hc4944aa7, 32'h43b1d5a4} /* (13, 30, 30) {real, imag} */,
  {32'hc1d7f900, 32'h42c4c2f2} /* (13, 30, 29) {real, imag} */,
  {32'h4326cde5, 32'hc2b97aac} /* (13, 30, 28) {real, imag} */,
  {32'hc34110e9, 32'hc2ebc80c} /* (13, 30, 27) {real, imag} */,
  {32'h42026cf1, 32'hc11628d0} /* (13, 30, 26) {real, imag} */,
  {32'h41aec43e, 32'hc1d381d0} /* (13, 30, 25) {real, imag} */,
  {32'hc28599e0, 32'h429c9582} /* (13, 30, 24) {real, imag} */,
  {32'hc24de024, 32'hc03f6a50} /* (13, 30, 23) {real, imag} */,
  {32'h42cfd1a5, 32'hc31b9266} /* (13, 30, 22) {real, imag} */,
  {32'hbfe328c0, 32'h417308fc} /* (13, 30, 21) {real, imag} */,
  {32'hc20fb1f8, 32'h432aec93} /* (13, 30, 20) {real, imag} */,
  {32'hc21d69d8, 32'hc276ad62} /* (13, 30, 19) {real, imag} */,
  {32'hc1bde2a3, 32'hc2263deb} /* (13, 30, 18) {real, imag} */,
  {32'hc084283c, 32'hc22ec59e} /* (13, 30, 17) {real, imag} */,
  {32'h4115d758, 32'h00000000} /* (13, 30, 16) {real, imag} */,
  {32'hc084283c, 32'h422ec59e} /* (13, 30, 15) {real, imag} */,
  {32'hc1bde2a3, 32'h42263deb} /* (13, 30, 14) {real, imag} */,
  {32'hc21d69d8, 32'h4276ad62} /* (13, 30, 13) {real, imag} */,
  {32'hc20fb1f8, 32'hc32aec93} /* (13, 30, 12) {real, imag} */,
  {32'hbfe328c0, 32'hc17308fc} /* (13, 30, 11) {real, imag} */,
  {32'h42cfd1a5, 32'h431b9266} /* (13, 30, 10) {real, imag} */,
  {32'hc24de024, 32'h403f6a50} /* (13, 30, 9) {real, imag} */,
  {32'hc28599e0, 32'hc29c9582} /* (13, 30, 8) {real, imag} */,
  {32'h41aec43e, 32'h41d381d0} /* (13, 30, 7) {real, imag} */,
  {32'h42026cf1, 32'h411628d0} /* (13, 30, 6) {real, imag} */,
  {32'hc34110e9, 32'h42ebc80c} /* (13, 30, 5) {real, imag} */,
  {32'h4326cde5, 32'h42b97aac} /* (13, 30, 4) {real, imag} */,
  {32'hc1d7f900, 32'hc2c4c2f2} /* (13, 30, 3) {real, imag} */,
  {32'hc4944aa7, 32'hc3b1d5a4} /* (13, 30, 2) {real, imag} */,
  {32'h4554571a, 32'h44abdc7e} /* (13, 30, 1) {real, imag} */,
  {32'h45789434, 32'h00000000} /* (13, 30, 0) {real, imag} */,
  {32'h45671dcf, 32'hc47f0678} /* (13, 29, 31) {real, imag} */,
  {32'hc4a04b8a, 32'h43a1fffe} /* (13, 29, 30) {real, imag} */,
  {32'h43258a0f, 32'h42d638ce} /* (13, 29, 29) {real, imag} */,
  {32'h431155ed, 32'hc29d3845} /* (13, 29, 28) {real, imag} */,
  {32'hc30dd511, 32'hc032f510} /* (13, 29, 27) {real, imag} */,
  {32'h40625bcc, 32'hc1f090ac} /* (13, 29, 26) {real, imag} */,
  {32'hc0295948, 32'hc205c89f} /* (13, 29, 25) {real, imag} */,
  {32'hc3554480, 32'h43298d62} /* (13, 29, 24) {real, imag} */,
  {32'hc2a3ff15, 32'h4302d5f7} /* (13, 29, 23) {real, imag} */,
  {32'h4242cacf, 32'hc13b9a5a} /* (13, 29, 22) {real, imag} */,
  {32'hc150c70a, 32'h41dcc9c8} /* (13, 29, 21) {real, imag} */,
  {32'hc2830fd2, 32'h4180add6} /* (13, 29, 20) {real, imag} */,
  {32'hc2a6f722, 32'hc143fb54} /* (13, 29, 19) {real, imag} */,
  {32'h41b22a4a, 32'hc24c5fb5} /* (13, 29, 18) {real, imag} */,
  {32'hc29e59d4, 32'hc1170ce2} /* (13, 29, 17) {real, imag} */,
  {32'hc20ba8f7, 32'h00000000} /* (13, 29, 16) {real, imag} */,
  {32'hc29e59d4, 32'h41170ce2} /* (13, 29, 15) {real, imag} */,
  {32'h41b22a4a, 32'h424c5fb5} /* (13, 29, 14) {real, imag} */,
  {32'hc2a6f722, 32'h4143fb54} /* (13, 29, 13) {real, imag} */,
  {32'hc2830fd2, 32'hc180add6} /* (13, 29, 12) {real, imag} */,
  {32'hc150c70a, 32'hc1dcc9c8} /* (13, 29, 11) {real, imag} */,
  {32'h4242cacf, 32'h413b9a5a} /* (13, 29, 10) {real, imag} */,
  {32'hc2a3ff15, 32'hc302d5f7} /* (13, 29, 9) {real, imag} */,
  {32'hc3554480, 32'hc3298d62} /* (13, 29, 8) {real, imag} */,
  {32'hc0295948, 32'h4205c89f} /* (13, 29, 7) {real, imag} */,
  {32'h40625bcc, 32'h41f090ac} /* (13, 29, 6) {real, imag} */,
  {32'hc30dd511, 32'h4032f510} /* (13, 29, 5) {real, imag} */,
  {32'h431155ed, 32'h429d3845} /* (13, 29, 4) {real, imag} */,
  {32'h43258a0f, 32'hc2d638ce} /* (13, 29, 3) {real, imag} */,
  {32'hc4a04b8a, 32'hc3a1fffe} /* (13, 29, 2) {real, imag} */,
  {32'h45671dcf, 32'h447f0678} /* (13, 29, 1) {real, imag} */,
  {32'h457c6bc2, 32'h00000000} /* (13, 29, 0) {real, imag} */,
  {32'h456d3b6c, 32'hc4638032} /* (13, 28, 31) {real, imag} */,
  {32'hc4aecae2, 32'h43826f26} /* (13, 28, 30) {real, imag} */,
  {32'hc08dc15c, 32'hc187b0f6} /* (13, 28, 29) {real, imag} */,
  {32'h42678c54, 32'hc34226f3} /* (13, 28, 28) {real, imag} */,
  {32'hc23351a6, 32'h4279e24c} /* (13, 28, 27) {real, imag} */,
  {32'h42295226, 32'h4132863c} /* (13, 28, 26) {real, imag} */,
  {32'h42337aa7, 32'h4204a6ff} /* (13, 28, 25) {real, imag} */,
  {32'hc1f8c841, 32'h42f2c819} /* (13, 28, 24) {real, imag} */,
  {32'hc2d6c8c1, 32'h4035ce98} /* (13, 28, 23) {real, imag} */,
  {32'hc2d30a0e, 32'h41a35150} /* (13, 28, 22) {real, imag} */,
  {32'hc1808339, 32'h40816bc8} /* (13, 28, 21) {real, imag} */,
  {32'h42264821, 32'hc29f1d6d} /* (13, 28, 20) {real, imag} */,
  {32'h4286bfa4, 32'hc1296497} /* (13, 28, 19) {real, imag} */,
  {32'h420cfa14, 32'h426d6668} /* (13, 28, 18) {real, imag} */,
  {32'h4215c4e2, 32'h41a6fa94} /* (13, 28, 17) {real, imag} */,
  {32'hc256ce0a, 32'h00000000} /* (13, 28, 16) {real, imag} */,
  {32'h4215c4e2, 32'hc1a6fa94} /* (13, 28, 15) {real, imag} */,
  {32'h420cfa14, 32'hc26d6668} /* (13, 28, 14) {real, imag} */,
  {32'h4286bfa4, 32'h41296497} /* (13, 28, 13) {real, imag} */,
  {32'h42264821, 32'h429f1d6d} /* (13, 28, 12) {real, imag} */,
  {32'hc1808339, 32'hc0816bc8} /* (13, 28, 11) {real, imag} */,
  {32'hc2d30a0e, 32'hc1a35150} /* (13, 28, 10) {real, imag} */,
  {32'hc2d6c8c1, 32'hc035ce98} /* (13, 28, 9) {real, imag} */,
  {32'hc1f8c841, 32'hc2f2c819} /* (13, 28, 8) {real, imag} */,
  {32'h42337aa7, 32'hc204a6ff} /* (13, 28, 7) {real, imag} */,
  {32'h42295226, 32'hc132863c} /* (13, 28, 6) {real, imag} */,
  {32'hc23351a6, 32'hc279e24c} /* (13, 28, 5) {real, imag} */,
  {32'h42678c54, 32'h434226f3} /* (13, 28, 4) {real, imag} */,
  {32'hc08dc15c, 32'h4187b0f6} /* (13, 28, 3) {real, imag} */,
  {32'hc4aecae2, 32'hc3826f26} /* (13, 28, 2) {real, imag} */,
  {32'h456d3b6c, 32'h44638032} /* (13, 28, 1) {real, imag} */,
  {32'h4574286a, 32'h00000000} /* (13, 28, 0) {real, imag} */,
  {32'h457069b0, 32'hc45d5c91} /* (13, 27, 31) {real, imag} */,
  {32'hc4bbdd31, 32'h434e3804} /* (13, 27, 30) {real, imag} */,
  {32'h41bca0c0, 32'hc3025356} /* (13, 27, 29) {real, imag} */,
  {32'h42588a80, 32'hc3375fa6} /* (13, 27, 28) {real, imag} */,
  {32'hc2f25d0a, 32'h432e7522} /* (13, 27, 27) {real, imag} */,
  {32'hc233f0c4, 32'h4225a00b} /* (13, 27, 26) {real, imag} */,
  {32'h42ae90b4, 32'hc1da6f8a} /* (13, 27, 25) {real, imag} */,
  {32'h419e0cde, 32'h426d2dd7} /* (13, 27, 24) {real, imag} */,
  {32'h419ea78e, 32'hc2b5d36b} /* (13, 27, 23) {real, imag} */,
  {32'h42c533da, 32'hc1370094} /* (13, 27, 22) {real, imag} */,
  {32'hc2a6fa04, 32'h4209470c} /* (13, 27, 21) {real, imag} */,
  {32'h42a54166, 32'h4318f85e} /* (13, 27, 20) {real, imag} */,
  {32'h422a8f18, 32'hc142d820} /* (13, 27, 19) {real, imag} */,
  {32'h424dbd5f, 32'h41256713} /* (13, 27, 18) {real, imag} */,
  {32'hc2a29b71, 32'h40048c68} /* (13, 27, 17) {real, imag} */,
  {32'h4226d8b2, 32'h00000000} /* (13, 27, 16) {real, imag} */,
  {32'hc2a29b71, 32'hc0048c68} /* (13, 27, 15) {real, imag} */,
  {32'h424dbd5f, 32'hc1256713} /* (13, 27, 14) {real, imag} */,
  {32'h422a8f18, 32'h4142d820} /* (13, 27, 13) {real, imag} */,
  {32'h42a54166, 32'hc318f85e} /* (13, 27, 12) {real, imag} */,
  {32'hc2a6fa04, 32'hc209470c} /* (13, 27, 11) {real, imag} */,
  {32'h42c533da, 32'h41370094} /* (13, 27, 10) {real, imag} */,
  {32'h419ea78e, 32'h42b5d36b} /* (13, 27, 9) {real, imag} */,
  {32'h419e0cde, 32'hc26d2dd7} /* (13, 27, 8) {real, imag} */,
  {32'h42ae90b4, 32'h41da6f8a} /* (13, 27, 7) {real, imag} */,
  {32'hc233f0c4, 32'hc225a00b} /* (13, 27, 6) {real, imag} */,
  {32'hc2f25d0a, 32'hc32e7522} /* (13, 27, 5) {real, imag} */,
  {32'h42588a80, 32'h43375fa6} /* (13, 27, 4) {real, imag} */,
  {32'h41bca0c0, 32'h43025356} /* (13, 27, 3) {real, imag} */,
  {32'hc4bbdd31, 32'hc34e3804} /* (13, 27, 2) {real, imag} */,
  {32'h457069b0, 32'h445d5c91} /* (13, 27, 1) {real, imag} */,
  {32'h45760581, 32'h00000000} /* (13, 27, 0) {real, imag} */,
  {32'h456fb89a, 32'hc4307fa5} /* (13, 26, 31) {real, imag} */,
  {32'hc4c6962a, 32'h4333078e} /* (13, 26, 30) {real, imag} */,
  {32'hc2ace63a, 32'hc293c3c6} /* (13, 26, 29) {real, imag} */,
  {32'h43056ad7, 32'hc33ec25f} /* (13, 26, 28) {real, imag} */,
  {32'hc2756067, 32'h42eff9be} /* (13, 26, 27) {real, imag} */,
  {32'hc2bddc62, 32'hc2308716} /* (13, 26, 26) {real, imag} */,
  {32'hc207b8f0, 32'hc24e71bb} /* (13, 26, 25) {real, imag} */,
  {32'hc3263c5e, 32'h42ae3535} /* (13, 26, 24) {real, imag} */,
  {32'h4201e583, 32'h428938da} /* (13, 26, 23) {real, imag} */,
  {32'h429cfda6, 32'h428d87e3} /* (13, 26, 22) {real, imag} */,
  {32'hc29b5c22, 32'hc34750b4} /* (13, 26, 21) {real, imag} */,
  {32'hc2536dc8, 32'h4175fa96} /* (13, 26, 20) {real, imag} */,
  {32'hc0927834, 32'h4140eeb8} /* (13, 26, 19) {real, imag} */,
  {32'h4199e129, 32'hc11cc34a} /* (13, 26, 18) {real, imag} */,
  {32'h4200b408, 32'h41f444bb} /* (13, 26, 17) {real, imag} */,
  {32'hc29886fa, 32'h00000000} /* (13, 26, 16) {real, imag} */,
  {32'h4200b408, 32'hc1f444bb} /* (13, 26, 15) {real, imag} */,
  {32'h4199e129, 32'h411cc34a} /* (13, 26, 14) {real, imag} */,
  {32'hc0927834, 32'hc140eeb8} /* (13, 26, 13) {real, imag} */,
  {32'hc2536dc8, 32'hc175fa96} /* (13, 26, 12) {real, imag} */,
  {32'hc29b5c22, 32'h434750b4} /* (13, 26, 11) {real, imag} */,
  {32'h429cfda6, 32'hc28d87e3} /* (13, 26, 10) {real, imag} */,
  {32'h4201e583, 32'hc28938da} /* (13, 26, 9) {real, imag} */,
  {32'hc3263c5e, 32'hc2ae3535} /* (13, 26, 8) {real, imag} */,
  {32'hc207b8f0, 32'h424e71bb} /* (13, 26, 7) {real, imag} */,
  {32'hc2bddc62, 32'h42308716} /* (13, 26, 6) {real, imag} */,
  {32'hc2756067, 32'hc2eff9be} /* (13, 26, 5) {real, imag} */,
  {32'h43056ad7, 32'h433ec25f} /* (13, 26, 4) {real, imag} */,
  {32'hc2ace63a, 32'h4293c3c6} /* (13, 26, 3) {real, imag} */,
  {32'hc4c6962a, 32'hc333078e} /* (13, 26, 2) {real, imag} */,
  {32'h456fb89a, 32'h44307fa5} /* (13, 26, 1) {real, imag} */,
  {32'h4568a0c4, 32'h00000000} /* (13, 26, 0) {real, imag} */,
  {32'h4568c330, 32'hc42aee1b} /* (13, 25, 31) {real, imag} */,
  {32'hc4c36562, 32'h43748719} /* (13, 25, 30) {real, imag} */,
  {32'hc24880fe, 32'hc2e349e0} /* (13, 25, 29) {real, imag} */,
  {32'h436c7139, 32'hc2df8180} /* (13, 25, 28) {real, imag} */,
  {32'hc34bce94, 32'h42b25794} /* (13, 25, 27) {real, imag} */,
  {32'hc1e83300, 32'hc2f3ad08} /* (13, 25, 26) {real, imag} */,
  {32'h4148a408, 32'hc184c29c} /* (13, 25, 25) {real, imag} */,
  {32'hc0e80850, 32'h43015cfb} /* (13, 25, 24) {real, imag} */,
  {32'h4299563a, 32'h42d39d42} /* (13, 25, 23) {real, imag} */,
  {32'hc2bd6f96, 32'hc27798a3} /* (13, 25, 22) {real, imag} */,
  {32'h429f039a, 32'hc194f9b0} /* (13, 25, 21) {real, imag} */,
  {32'h411f037a, 32'h40a5ae58} /* (13, 25, 20) {real, imag} */,
  {32'h4241c991, 32'hc206889a} /* (13, 25, 19) {real, imag} */,
  {32'hbf67db60, 32'h42495192} /* (13, 25, 18) {real, imag} */,
  {32'hc28d7883, 32'hc28bc598} /* (13, 25, 17) {real, imag} */,
  {32'hc291057a, 32'h00000000} /* (13, 25, 16) {real, imag} */,
  {32'hc28d7883, 32'h428bc598} /* (13, 25, 15) {real, imag} */,
  {32'hbf67db60, 32'hc2495192} /* (13, 25, 14) {real, imag} */,
  {32'h4241c991, 32'h4206889a} /* (13, 25, 13) {real, imag} */,
  {32'h411f037a, 32'hc0a5ae58} /* (13, 25, 12) {real, imag} */,
  {32'h429f039a, 32'h4194f9b0} /* (13, 25, 11) {real, imag} */,
  {32'hc2bd6f96, 32'h427798a3} /* (13, 25, 10) {real, imag} */,
  {32'h4299563a, 32'hc2d39d42} /* (13, 25, 9) {real, imag} */,
  {32'hc0e80850, 32'hc3015cfb} /* (13, 25, 8) {real, imag} */,
  {32'h4148a408, 32'h4184c29c} /* (13, 25, 7) {real, imag} */,
  {32'hc1e83300, 32'h42f3ad08} /* (13, 25, 6) {real, imag} */,
  {32'hc34bce94, 32'hc2b25794} /* (13, 25, 5) {real, imag} */,
  {32'h436c7139, 32'h42df8180} /* (13, 25, 4) {real, imag} */,
  {32'hc24880fe, 32'h42e349e0} /* (13, 25, 3) {real, imag} */,
  {32'hc4c36562, 32'hc3748719} /* (13, 25, 2) {real, imag} */,
  {32'h4568c330, 32'h442aee1b} /* (13, 25, 1) {real, imag} */,
  {32'h455378e4, 32'h00000000} /* (13, 25, 0) {real, imag} */,
  {32'h4554d23d, 32'hc42b1978} /* (13, 24, 31) {real, imag} */,
  {32'hc4bc5d71, 32'h43b74457} /* (13, 24, 30) {real, imag} */,
  {32'h417abfec, 32'hc356ca8e} /* (13, 24, 29) {real, imag} */,
  {32'h43849e7c, 32'hc28dac74} /* (13, 24, 28) {real, imag} */,
  {32'hc362045e, 32'h432c8c35} /* (13, 24, 27) {real, imag} */,
  {32'hc2326f5f, 32'hc34bed18} /* (13, 24, 26) {real, imag} */,
  {32'h4242e1db, 32'h4296f9e1} /* (13, 24, 25) {real, imag} */,
  {32'h42125b14, 32'h427a24ee} /* (13, 24, 24) {real, imag} */,
  {32'h431ef564, 32'h421c0cc4} /* (13, 24, 23) {real, imag} */,
  {32'hc26d0132, 32'hc21b975d} /* (13, 24, 22) {real, imag} */,
  {32'h426e6cea, 32'h4228e994} /* (13, 24, 21) {real, imag} */,
  {32'hc2097840, 32'h4163a864} /* (13, 24, 20) {real, imag} */,
  {32'h42158132, 32'hc2f9223e} /* (13, 24, 19) {real, imag} */,
  {32'hc223750c, 32'h4214b87e} /* (13, 24, 18) {real, imag} */,
  {32'hc00bf3e0, 32'h414942c2} /* (13, 24, 17) {real, imag} */,
  {32'h41e3f4ea, 32'h00000000} /* (13, 24, 16) {real, imag} */,
  {32'hc00bf3e0, 32'hc14942c2} /* (13, 24, 15) {real, imag} */,
  {32'hc223750c, 32'hc214b87e} /* (13, 24, 14) {real, imag} */,
  {32'h42158132, 32'h42f9223e} /* (13, 24, 13) {real, imag} */,
  {32'hc2097840, 32'hc163a864} /* (13, 24, 12) {real, imag} */,
  {32'h426e6cea, 32'hc228e994} /* (13, 24, 11) {real, imag} */,
  {32'hc26d0132, 32'h421b975d} /* (13, 24, 10) {real, imag} */,
  {32'h431ef564, 32'hc21c0cc4} /* (13, 24, 9) {real, imag} */,
  {32'h42125b14, 32'hc27a24ee} /* (13, 24, 8) {real, imag} */,
  {32'h4242e1db, 32'hc296f9e1} /* (13, 24, 7) {real, imag} */,
  {32'hc2326f5f, 32'h434bed18} /* (13, 24, 6) {real, imag} */,
  {32'hc362045e, 32'hc32c8c35} /* (13, 24, 5) {real, imag} */,
  {32'h43849e7c, 32'h428dac74} /* (13, 24, 4) {real, imag} */,
  {32'h417abfec, 32'h4356ca8e} /* (13, 24, 3) {real, imag} */,
  {32'hc4bc5d71, 32'hc3b74457} /* (13, 24, 2) {real, imag} */,
  {32'h4554d23d, 32'h442b1978} /* (13, 24, 1) {real, imag} */,
  {32'h45266250, 32'h00000000} /* (13, 24, 0) {real, imag} */,
  {32'h45320657, 32'hc3e5cbde} /* (13, 23, 31) {real, imag} */,
  {32'hc49083ed, 32'h43b9a7bc} /* (13, 23, 30) {real, imag} */,
  {32'hc283cba6, 32'hc3327d54} /* (13, 23, 29) {real, imag} */,
  {32'h438007d2, 32'hc315ef53} /* (13, 23, 28) {real, imag} */,
  {32'hc32639c9, 32'h42b59888} /* (13, 23, 27) {real, imag} */,
  {32'hc2ace850, 32'h407307f8} /* (13, 23, 26) {real, imag} */,
  {32'h41d68292, 32'hc2843a43} /* (13, 23, 25) {real, imag} */,
  {32'hc256b61b, 32'h41c1ab04} /* (13, 23, 24) {real, imag} */,
  {32'h421c0529, 32'h4243ce59} /* (13, 23, 23) {real, imag} */,
  {32'hc25dacd3, 32'h4195c762} /* (13, 23, 22) {real, imag} */,
  {32'hc22f048f, 32'h4103cab0} /* (13, 23, 21) {real, imag} */,
  {32'h424158a6, 32'h418b7bfa} /* (13, 23, 20) {real, imag} */,
  {32'hc211d11c, 32'h41a49524} /* (13, 23, 19) {real, imag} */,
  {32'hc13378b8, 32'h42c66907} /* (13, 23, 18) {real, imag} */,
  {32'h426814dc, 32'hc1d6ec17} /* (13, 23, 17) {real, imag} */,
  {32'h422ae316, 32'h00000000} /* (13, 23, 16) {real, imag} */,
  {32'h426814dc, 32'h41d6ec17} /* (13, 23, 15) {real, imag} */,
  {32'hc13378b8, 32'hc2c66907} /* (13, 23, 14) {real, imag} */,
  {32'hc211d11c, 32'hc1a49524} /* (13, 23, 13) {real, imag} */,
  {32'h424158a6, 32'hc18b7bfa} /* (13, 23, 12) {real, imag} */,
  {32'hc22f048f, 32'hc103cab0} /* (13, 23, 11) {real, imag} */,
  {32'hc25dacd3, 32'hc195c762} /* (13, 23, 10) {real, imag} */,
  {32'h421c0529, 32'hc243ce59} /* (13, 23, 9) {real, imag} */,
  {32'hc256b61b, 32'hc1c1ab04} /* (13, 23, 8) {real, imag} */,
  {32'h41d68292, 32'h42843a43} /* (13, 23, 7) {real, imag} */,
  {32'hc2ace850, 32'hc07307f8} /* (13, 23, 6) {real, imag} */,
  {32'hc32639c9, 32'hc2b59888} /* (13, 23, 5) {real, imag} */,
  {32'h438007d2, 32'h4315ef53} /* (13, 23, 4) {real, imag} */,
  {32'hc283cba6, 32'h43327d54} /* (13, 23, 3) {real, imag} */,
  {32'hc49083ed, 32'hc3b9a7bc} /* (13, 23, 2) {real, imag} */,
  {32'h45320657, 32'h43e5cbde} /* (13, 23, 1) {real, imag} */,
  {32'h4502e690, 32'h00000000} /* (13, 23, 0) {real, imag} */,
  {32'h44f6c0ec, 32'hc3811890} /* (13, 22, 31) {real, imag} */,
  {32'hc4317d09, 32'h431eb5ca} /* (13, 22, 30) {real, imag} */,
  {32'hc3008c1f, 32'hc2eef69c} /* (13, 22, 29) {real, imag} */,
  {32'h4377b5eb, 32'hc3755a27} /* (13, 22, 28) {real, imag} */,
  {32'hc354683b, 32'h42ec3032} /* (13, 22, 27) {real, imag} */,
  {32'hc29e26ea, 32'h424ec6cc} /* (13, 22, 26) {real, imag} */,
  {32'h404357e8, 32'hc1e58824} /* (13, 22, 25) {real, imag} */,
  {32'hc2b24034, 32'h4168b7c0} /* (13, 22, 24) {real, imag} */,
  {32'hc200df10, 32'h41bc50f0} /* (13, 22, 23) {real, imag} */,
  {32'h3ff4edd0, 32'hc26e44d4} /* (13, 22, 22) {real, imag} */,
  {32'hc2695f02, 32'h400cbc30} /* (13, 22, 21) {real, imag} */,
  {32'hc274e2cc, 32'hc1c1e116} /* (13, 22, 20) {real, imag} */,
  {32'hc25185c8, 32'hc2bb204a} /* (13, 22, 19) {real, imag} */,
  {32'h4216c0e6, 32'h4213f586} /* (13, 22, 18) {real, imag} */,
  {32'h42070778, 32'h4285d717} /* (13, 22, 17) {real, imag} */,
  {32'hc15bd7e6, 32'h00000000} /* (13, 22, 16) {real, imag} */,
  {32'h42070778, 32'hc285d717} /* (13, 22, 15) {real, imag} */,
  {32'h4216c0e6, 32'hc213f586} /* (13, 22, 14) {real, imag} */,
  {32'hc25185c8, 32'h42bb204a} /* (13, 22, 13) {real, imag} */,
  {32'hc274e2cc, 32'h41c1e116} /* (13, 22, 12) {real, imag} */,
  {32'hc2695f02, 32'hc00cbc30} /* (13, 22, 11) {real, imag} */,
  {32'h3ff4edd0, 32'h426e44d4} /* (13, 22, 10) {real, imag} */,
  {32'hc200df10, 32'hc1bc50f0} /* (13, 22, 9) {real, imag} */,
  {32'hc2b24034, 32'hc168b7c0} /* (13, 22, 8) {real, imag} */,
  {32'h404357e8, 32'h41e58824} /* (13, 22, 7) {real, imag} */,
  {32'hc29e26ea, 32'hc24ec6cc} /* (13, 22, 6) {real, imag} */,
  {32'hc354683b, 32'hc2ec3032} /* (13, 22, 5) {real, imag} */,
  {32'h4377b5eb, 32'h43755a27} /* (13, 22, 4) {real, imag} */,
  {32'hc3008c1f, 32'h42eef69c} /* (13, 22, 3) {real, imag} */,
  {32'hc4317d09, 32'hc31eb5ca} /* (13, 22, 2) {real, imag} */,
  {32'h44f6c0ec, 32'h43811890} /* (13, 22, 1) {real, imag} */,
  {32'h44bf6c7d, 32'h00000000} /* (13, 22, 0) {real, imag} */,
  {32'h4400e193, 32'h4214c690} /* (13, 21, 31) {real, imag} */,
  {32'hc34c8ffa, 32'h429c0b56} /* (13, 21, 30) {real, imag} */,
  {32'h4280f310, 32'hc2929b34} /* (13, 21, 29) {real, imag} */,
  {32'h43070504, 32'hc3081042} /* (13, 21, 28) {real, imag} */,
  {32'hc2b6e35e, 32'h431ebc2e} /* (13, 21, 27) {real, imag} */,
  {32'hc3011425, 32'hc1f7c973} /* (13, 21, 26) {real, imag} */,
  {32'h429f8a1d, 32'hc2840796} /* (13, 21, 25) {real, imag} */,
  {32'h432dddf4, 32'h4201fd1f} /* (13, 21, 24) {real, imag} */,
  {32'hc2a794de, 32'h423d7e70} /* (13, 21, 23) {real, imag} */,
  {32'hc2256dc2, 32'h421e84f7} /* (13, 21, 22) {real, imag} */,
  {32'h41fa1087, 32'h421193f4} /* (13, 21, 21) {real, imag} */,
  {32'h41d812a2, 32'hc280beeb} /* (13, 21, 20) {real, imag} */,
  {32'h42874389, 32'hc2aaf772} /* (13, 21, 19) {real, imag} */,
  {32'h418d453c, 32'hc211c38f} /* (13, 21, 18) {real, imag} */,
  {32'hc1f50bf5, 32'h42e4e644} /* (13, 21, 17) {real, imag} */,
  {32'h42771ea2, 32'h00000000} /* (13, 21, 16) {real, imag} */,
  {32'hc1f50bf5, 32'hc2e4e644} /* (13, 21, 15) {real, imag} */,
  {32'h418d453c, 32'h4211c38f} /* (13, 21, 14) {real, imag} */,
  {32'h42874389, 32'h42aaf772} /* (13, 21, 13) {real, imag} */,
  {32'h41d812a2, 32'h4280beeb} /* (13, 21, 12) {real, imag} */,
  {32'h41fa1087, 32'hc21193f4} /* (13, 21, 11) {real, imag} */,
  {32'hc2256dc2, 32'hc21e84f7} /* (13, 21, 10) {real, imag} */,
  {32'hc2a794de, 32'hc23d7e70} /* (13, 21, 9) {real, imag} */,
  {32'h432dddf4, 32'hc201fd1f} /* (13, 21, 8) {real, imag} */,
  {32'h429f8a1d, 32'h42840796} /* (13, 21, 7) {real, imag} */,
  {32'hc3011425, 32'h41f7c973} /* (13, 21, 6) {real, imag} */,
  {32'hc2b6e35e, 32'hc31ebc2e} /* (13, 21, 5) {real, imag} */,
  {32'h43070504, 32'h43081042} /* (13, 21, 4) {real, imag} */,
  {32'h4280f310, 32'h42929b34} /* (13, 21, 3) {real, imag} */,
  {32'hc34c8ffa, 32'hc29c0b56} /* (13, 21, 2) {real, imag} */,
  {32'h4400e193, 32'hc214c690} /* (13, 21, 1) {real, imag} */,
  {32'h441c3f21, 32'h00000000} /* (13, 21, 0) {real, imag} */,
  {32'hc4966038, 32'h431eabec} /* (13, 20, 31) {real, imag} */,
  {32'h43faf4d0, 32'hc2c64c9a} /* (13, 20, 30) {real, imag} */,
  {32'h42529b22, 32'hc259efb3} /* (13, 20, 29) {real, imag} */,
  {32'h41d3bf44, 32'h4151e390} /* (13, 20, 28) {real, imag} */,
  {32'h42f31331, 32'hc2ec32d0} /* (13, 20, 27) {real, imag} */,
  {32'hc2c617d4, 32'hc236dcd9} /* (13, 20, 26) {real, imag} */,
  {32'h41a90b80, 32'hc25a1db7} /* (13, 20, 25) {real, imag} */,
  {32'h42820d34, 32'hc180045c} /* (13, 20, 24) {real, imag} */,
  {32'h419fe4c1, 32'h4203d9a6} /* (13, 20, 23) {real, imag} */,
  {32'hc216da4e, 32'h4186eab4} /* (13, 20, 22) {real, imag} */,
  {32'h42fc40b8, 32'h3f616b60} /* (13, 20, 21) {real, imag} */,
  {32'h4139733d, 32'h4266e60f} /* (13, 20, 20) {real, imag} */,
  {32'hc2380564, 32'hc20bac25} /* (13, 20, 19) {real, imag} */,
  {32'h416dda82, 32'h41644472} /* (13, 20, 18) {real, imag} */,
  {32'hc27ced3b, 32'h42725aff} /* (13, 20, 17) {real, imag} */,
  {32'hc2513a42, 32'h00000000} /* (13, 20, 16) {real, imag} */,
  {32'hc27ced3b, 32'hc2725aff} /* (13, 20, 15) {real, imag} */,
  {32'h416dda82, 32'hc1644472} /* (13, 20, 14) {real, imag} */,
  {32'hc2380564, 32'h420bac25} /* (13, 20, 13) {real, imag} */,
  {32'h4139733d, 32'hc266e60f} /* (13, 20, 12) {real, imag} */,
  {32'h42fc40b8, 32'hbf616b60} /* (13, 20, 11) {real, imag} */,
  {32'hc216da4e, 32'hc186eab4} /* (13, 20, 10) {real, imag} */,
  {32'h419fe4c1, 32'hc203d9a6} /* (13, 20, 9) {real, imag} */,
  {32'h42820d34, 32'h4180045c} /* (13, 20, 8) {real, imag} */,
  {32'h41a90b80, 32'h425a1db7} /* (13, 20, 7) {real, imag} */,
  {32'hc2c617d4, 32'h4236dcd9} /* (13, 20, 6) {real, imag} */,
  {32'h42f31331, 32'h42ec32d0} /* (13, 20, 5) {real, imag} */,
  {32'h41d3bf44, 32'hc151e390} /* (13, 20, 4) {real, imag} */,
  {32'h42529b22, 32'h4259efb3} /* (13, 20, 3) {real, imag} */,
  {32'h43faf4d0, 32'h42c64c9a} /* (13, 20, 2) {real, imag} */,
  {32'hc4966038, 32'hc31eabec} /* (13, 20, 1) {real, imag} */,
  {32'hc433eae2, 32'h00000000} /* (13, 20, 0) {real, imag} */,
  {32'hc5065280, 32'h438e7cc2} /* (13, 19, 31) {real, imag} */,
  {32'h4471bcd4, 32'hc30ed1c3} /* (13, 19, 30) {real, imag} */,
  {32'h420054a8, 32'hc133cbec} /* (13, 19, 29) {real, imag} */,
  {32'hc2935e99, 32'h4316cdaf} /* (13, 19, 28) {real, imag} */,
  {32'h435b5159, 32'hc32d488a} /* (13, 19, 27) {real, imag} */,
  {32'h4140f5a6, 32'hc3062c89} /* (13, 19, 26) {real, imag} */,
  {32'h40a509e4, 32'h41d02ab2} /* (13, 19, 25) {real, imag} */,
  {32'h424d7931, 32'hc29793a8} /* (13, 19, 24) {real, imag} */,
  {32'h40828e38, 32'h42e49cb8} /* (13, 19, 23) {real, imag} */,
  {32'hc24c6bac, 32'hc2bd0a7f} /* (13, 19, 22) {real, imag} */,
  {32'h4236d62a, 32'hc11485c0} /* (13, 19, 21) {real, imag} */,
  {32'hc213279e, 32'h42a3918e} /* (13, 19, 20) {real, imag} */,
  {32'hc2766db6, 32'h418be880} /* (13, 19, 19) {real, imag} */,
  {32'hc205dc3d, 32'h4183dd92} /* (13, 19, 18) {real, imag} */,
  {32'h4184f8de, 32'hc0a17b54} /* (13, 19, 17) {real, imag} */,
  {32'h42f0c498, 32'h00000000} /* (13, 19, 16) {real, imag} */,
  {32'h4184f8de, 32'h40a17b54} /* (13, 19, 15) {real, imag} */,
  {32'hc205dc3d, 32'hc183dd92} /* (13, 19, 14) {real, imag} */,
  {32'hc2766db6, 32'hc18be880} /* (13, 19, 13) {real, imag} */,
  {32'hc213279e, 32'hc2a3918e} /* (13, 19, 12) {real, imag} */,
  {32'h4236d62a, 32'h411485c0} /* (13, 19, 11) {real, imag} */,
  {32'hc24c6bac, 32'h42bd0a7f} /* (13, 19, 10) {real, imag} */,
  {32'h40828e38, 32'hc2e49cb8} /* (13, 19, 9) {real, imag} */,
  {32'h424d7931, 32'h429793a8} /* (13, 19, 8) {real, imag} */,
  {32'h40a509e4, 32'hc1d02ab2} /* (13, 19, 7) {real, imag} */,
  {32'h4140f5a6, 32'h43062c89} /* (13, 19, 6) {real, imag} */,
  {32'h435b5159, 32'h432d488a} /* (13, 19, 5) {real, imag} */,
  {32'hc2935e99, 32'hc316cdaf} /* (13, 19, 4) {real, imag} */,
  {32'h420054a8, 32'h4133cbec} /* (13, 19, 3) {real, imag} */,
  {32'h4471bcd4, 32'h430ed1c3} /* (13, 19, 2) {real, imag} */,
  {32'hc5065280, 32'hc38e7cc2} /* (13, 19, 1) {real, imag} */,
  {32'hc4b4d430, 32'h00000000} /* (13, 19, 0) {real, imag} */,
  {32'hc528d5da, 32'h43b9f0f8} /* (13, 18, 31) {real, imag} */,
  {32'h44964f49, 32'hc3acde47} /* (13, 18, 30) {real, imag} */,
  {32'h42c31369, 32'hc28218d4} /* (13, 18, 29) {real, imag} */,
  {32'hc3133b25, 32'h432f01a8} /* (13, 18, 28) {real, imag} */,
  {32'h436b1034, 32'hc223afa3} /* (13, 18, 27) {real, imag} */,
  {32'h41189864, 32'hc1ead3a8} /* (13, 18, 26) {real, imag} */,
  {32'hc2635674, 32'h41c2ddd2} /* (13, 18, 25) {real, imag} */,
  {32'h42357f70, 32'hc29a3967} /* (13, 18, 24) {real, imag} */,
  {32'h426a2e8c, 32'hc08173ae} /* (13, 18, 23) {real, imag} */,
  {32'h42a37dca, 32'hc0e86d50} /* (13, 18, 22) {real, imag} */,
  {32'hc27d0868, 32'hc28ab974} /* (13, 18, 21) {real, imag} */,
  {32'h411c9acc, 32'h428fef06} /* (13, 18, 20) {real, imag} */,
  {32'hc26bfffc, 32'hc24795d8} /* (13, 18, 19) {real, imag} */,
  {32'h41a724a3, 32'hc260189a} /* (13, 18, 18) {real, imag} */,
  {32'hc1932242, 32'h42188ef3} /* (13, 18, 17) {real, imag} */,
  {32'hc2c6ed9e, 32'h00000000} /* (13, 18, 16) {real, imag} */,
  {32'hc1932242, 32'hc2188ef3} /* (13, 18, 15) {real, imag} */,
  {32'h41a724a3, 32'h4260189a} /* (13, 18, 14) {real, imag} */,
  {32'hc26bfffc, 32'h424795d8} /* (13, 18, 13) {real, imag} */,
  {32'h411c9acc, 32'hc28fef06} /* (13, 18, 12) {real, imag} */,
  {32'hc27d0868, 32'h428ab974} /* (13, 18, 11) {real, imag} */,
  {32'h42a37dca, 32'h40e86d50} /* (13, 18, 10) {real, imag} */,
  {32'h426a2e8c, 32'h408173ae} /* (13, 18, 9) {real, imag} */,
  {32'h42357f70, 32'h429a3967} /* (13, 18, 8) {real, imag} */,
  {32'hc2635674, 32'hc1c2ddd2} /* (13, 18, 7) {real, imag} */,
  {32'h41189864, 32'h41ead3a8} /* (13, 18, 6) {real, imag} */,
  {32'h436b1034, 32'h4223afa3} /* (13, 18, 5) {real, imag} */,
  {32'hc3133b25, 32'hc32f01a8} /* (13, 18, 4) {real, imag} */,
  {32'h42c31369, 32'h428218d4} /* (13, 18, 3) {real, imag} */,
  {32'h44964f49, 32'h43acde47} /* (13, 18, 2) {real, imag} */,
  {32'hc528d5da, 32'hc3b9f0f8} /* (13, 18, 1) {real, imag} */,
  {32'hc50392bc, 32'h00000000} /* (13, 18, 0) {real, imag} */,
  {32'hc542bccb, 32'h43d1b05e} /* (13, 17, 31) {real, imag} */,
  {32'h44ad2e9e, 32'hc3a89e34} /* (13, 17, 30) {real, imag} */,
  {32'h42e91d5e, 32'hc27a0d72} /* (13, 17, 29) {real, imag} */,
  {32'hc3169be6, 32'h4378a459} /* (13, 17, 28) {real, imag} */,
  {32'h43659f9e, 32'hc21c2f5e} /* (13, 17, 27) {real, imag} */,
  {32'h426efcc4, 32'hc2d778cf} /* (13, 17, 26) {real, imag} */,
  {32'hc2f66f89, 32'h41b268d3} /* (13, 17, 25) {real, imag} */,
  {32'h42a56258, 32'hc27ef44c} /* (13, 17, 24) {real, imag} */,
  {32'h41c3d3a4, 32'hc24b55e5} /* (13, 17, 23) {real, imag} */,
  {32'hc29fbdeb, 32'hc2a40ba8} /* (13, 17, 22) {real, imag} */,
  {32'hc28b866c, 32'hc25c348f} /* (13, 17, 21) {real, imag} */,
  {32'hc252bea0, 32'hc25e7f54} /* (13, 17, 20) {real, imag} */,
  {32'h41c8da66, 32'hbeb0d9c0} /* (13, 17, 19) {real, imag} */,
  {32'h42fdca50, 32'h42e9cb1b} /* (13, 17, 18) {real, imag} */,
  {32'h42965c44, 32'hc1785234} /* (13, 17, 17) {real, imag} */,
  {32'hc289af40, 32'h00000000} /* (13, 17, 16) {real, imag} */,
  {32'h42965c44, 32'h41785234} /* (13, 17, 15) {real, imag} */,
  {32'h42fdca50, 32'hc2e9cb1b} /* (13, 17, 14) {real, imag} */,
  {32'h41c8da66, 32'h3eb0d9c0} /* (13, 17, 13) {real, imag} */,
  {32'hc252bea0, 32'h425e7f54} /* (13, 17, 12) {real, imag} */,
  {32'hc28b866c, 32'h425c348f} /* (13, 17, 11) {real, imag} */,
  {32'hc29fbdeb, 32'h42a40ba8} /* (13, 17, 10) {real, imag} */,
  {32'h41c3d3a4, 32'h424b55e5} /* (13, 17, 9) {real, imag} */,
  {32'h42a56258, 32'h427ef44c} /* (13, 17, 8) {real, imag} */,
  {32'hc2f66f89, 32'hc1b268d3} /* (13, 17, 7) {real, imag} */,
  {32'h426efcc4, 32'h42d778cf} /* (13, 17, 6) {real, imag} */,
  {32'h43659f9e, 32'h421c2f5e} /* (13, 17, 5) {real, imag} */,
  {32'hc3169be6, 32'hc378a459} /* (13, 17, 4) {real, imag} */,
  {32'h42e91d5e, 32'h427a0d72} /* (13, 17, 3) {real, imag} */,
  {32'h44ad2e9e, 32'h43a89e34} /* (13, 17, 2) {real, imag} */,
  {32'hc542bccb, 32'hc3d1b05e} /* (13, 17, 1) {real, imag} */,
  {32'hc5231140, 32'h00000000} /* (13, 17, 0) {real, imag} */,
  {32'hc5571582, 32'h44132e0a} /* (13, 16, 31) {real, imag} */,
  {32'h44b0a2e2, 32'hc38bd41a} /* (13, 16, 30) {real, imag} */,
  {32'h42aa4e0b, 32'hc300dec2} /* (13, 16, 29) {real, imag} */,
  {32'hc32634ed, 32'h433d9ad6} /* (13, 16, 28) {real, imag} */,
  {32'h43053d12, 32'hc2e11dbe} /* (13, 16, 27) {real, imag} */,
  {32'h4218473c, 32'hc2930017} /* (13, 16, 26) {real, imag} */,
  {32'hc32e64d8, 32'h40bd00d8} /* (13, 16, 25) {real, imag} */,
  {32'h431669ae, 32'hc26244a9} /* (13, 16, 24) {real, imag} */,
  {32'hc0457690, 32'hc235b6d2} /* (13, 16, 23) {real, imag} */,
  {32'hc212b0c3, 32'h41d06a02} /* (13, 16, 22) {real, imag} */,
  {32'h42b0372b, 32'hc0d7fd94} /* (13, 16, 21) {real, imag} */,
  {32'hc2c48528, 32'hc29009e8} /* (13, 16, 20) {real, imag} */,
  {32'h42140281, 32'h41bcb255} /* (13, 16, 19) {real, imag} */,
  {32'hc18f5cf4, 32'h41d752b4} /* (13, 16, 18) {real, imag} */,
  {32'h42372db8, 32'hc2998222} /* (13, 16, 17) {real, imag} */,
  {32'h42082bce, 32'h00000000} /* (13, 16, 16) {real, imag} */,
  {32'h42372db8, 32'h42998222} /* (13, 16, 15) {real, imag} */,
  {32'hc18f5cf4, 32'hc1d752b4} /* (13, 16, 14) {real, imag} */,
  {32'h42140281, 32'hc1bcb255} /* (13, 16, 13) {real, imag} */,
  {32'hc2c48528, 32'h429009e8} /* (13, 16, 12) {real, imag} */,
  {32'h42b0372b, 32'h40d7fd94} /* (13, 16, 11) {real, imag} */,
  {32'hc212b0c3, 32'hc1d06a02} /* (13, 16, 10) {real, imag} */,
  {32'hc0457690, 32'h4235b6d2} /* (13, 16, 9) {real, imag} */,
  {32'h431669ae, 32'h426244a9} /* (13, 16, 8) {real, imag} */,
  {32'hc32e64d8, 32'hc0bd00d8} /* (13, 16, 7) {real, imag} */,
  {32'h4218473c, 32'h42930017} /* (13, 16, 6) {real, imag} */,
  {32'h43053d12, 32'h42e11dbe} /* (13, 16, 5) {real, imag} */,
  {32'hc32634ed, 32'hc33d9ad6} /* (13, 16, 4) {real, imag} */,
  {32'h42aa4e0b, 32'h4300dec2} /* (13, 16, 3) {real, imag} */,
  {32'h44b0a2e2, 32'h438bd41a} /* (13, 16, 2) {real, imag} */,
  {32'hc5571582, 32'hc4132e0a} /* (13, 16, 1) {real, imag} */,
  {32'hc519f5e5, 32'h00000000} /* (13, 16, 0) {real, imag} */,
  {32'hc5600e19, 32'h440145df} /* (13, 15, 31) {real, imag} */,
  {32'h449b6bf8, 32'hc36afe11} /* (13, 15, 30) {real, imag} */,
  {32'h418522e0, 32'h410efa58} /* (13, 15, 29) {real, imag} */,
  {32'hc34934a6, 32'h4360c6fb} /* (13, 15, 28) {real, imag} */,
  {32'h42ce1b44, 32'hc381ef06} /* (13, 15, 27) {real, imag} */,
  {32'hc1d27a20, 32'hc30c67d6} /* (13, 15, 26) {real, imag} */,
  {32'hc2aa65f1, 32'hc1c603cb} /* (13, 15, 25) {real, imag} */,
  {32'h42377113, 32'hc28fe7a2} /* (13, 15, 24) {real, imag} */,
  {32'hc1f295a8, 32'hc209bc63} /* (13, 15, 23) {real, imag} */,
  {32'hc2a18eab, 32'hbf3d7dc0} /* (13, 15, 22) {real, imag} */,
  {32'h4194fb46, 32'hc24ec647} /* (13, 15, 21) {real, imag} */,
  {32'h422f911a, 32'h40ceb640} /* (13, 15, 20) {real, imag} */,
  {32'h42daeeb2, 32'hc0da1e24} /* (13, 15, 19) {real, imag} */,
  {32'hc207d7a7, 32'h4124b348} /* (13, 15, 18) {real, imag} */,
  {32'h41c1cc18, 32'h426ea5cb} /* (13, 15, 17) {real, imag} */,
  {32'h42431d18, 32'h00000000} /* (13, 15, 16) {real, imag} */,
  {32'h41c1cc18, 32'hc26ea5cb} /* (13, 15, 15) {real, imag} */,
  {32'hc207d7a7, 32'hc124b348} /* (13, 15, 14) {real, imag} */,
  {32'h42daeeb2, 32'h40da1e24} /* (13, 15, 13) {real, imag} */,
  {32'h422f911a, 32'hc0ceb640} /* (13, 15, 12) {real, imag} */,
  {32'h4194fb46, 32'h424ec647} /* (13, 15, 11) {real, imag} */,
  {32'hc2a18eab, 32'h3f3d7dc0} /* (13, 15, 10) {real, imag} */,
  {32'hc1f295a8, 32'h4209bc63} /* (13, 15, 9) {real, imag} */,
  {32'h42377113, 32'h428fe7a2} /* (13, 15, 8) {real, imag} */,
  {32'hc2aa65f1, 32'h41c603cb} /* (13, 15, 7) {real, imag} */,
  {32'hc1d27a20, 32'h430c67d6} /* (13, 15, 6) {real, imag} */,
  {32'h42ce1b44, 32'h4381ef06} /* (13, 15, 5) {real, imag} */,
  {32'hc34934a6, 32'hc360c6fb} /* (13, 15, 4) {real, imag} */,
  {32'h418522e0, 32'hc10efa58} /* (13, 15, 3) {real, imag} */,
  {32'h449b6bf8, 32'h436afe11} /* (13, 15, 2) {real, imag} */,
  {32'hc5600e19, 32'hc40145df} /* (13, 15, 1) {real, imag} */,
  {32'hc5201d42, 32'h00000000} /* (13, 15, 0) {real, imag} */,
  {32'hc551ba7e, 32'h43813898} /* (13, 14, 31) {real, imag} */,
  {32'h44839641, 32'hc3457762} /* (13, 14, 30) {real, imag} */,
  {32'h413c3e48, 32'hc1e4a0ea} /* (13, 14, 29) {real, imag} */,
  {32'hc314b843, 32'h42807fd0} /* (13, 14, 28) {real, imag} */,
  {32'h42a6d26c, 32'hc2f14d76} /* (13, 14, 27) {real, imag} */,
  {32'h4034c520, 32'hc33bb03f} /* (13, 14, 26) {real, imag} */,
  {32'hc2facc9e, 32'hc2aacad4} /* (13, 14, 25) {real, imag} */,
  {32'h4057b9a0, 32'hc1c6fae8} /* (13, 14, 24) {real, imag} */,
  {32'hc220d328, 32'h41485a27} /* (13, 14, 23) {real, imag} */,
  {32'hc26dfe05, 32'hc297bd1d} /* (13, 14, 22) {real, imag} */,
  {32'hc2aa5e58, 32'h411a432c} /* (13, 14, 21) {real, imag} */,
  {32'h42c633ac, 32'hc1b8b4ec} /* (13, 14, 20) {real, imag} */,
  {32'hc283eff7, 32'hc1f7104c} /* (13, 14, 19) {real, imag} */,
  {32'hc0c02acc, 32'h40d97790} /* (13, 14, 18) {real, imag} */,
  {32'hc1a7668c, 32'h41d67262} /* (13, 14, 17) {real, imag} */,
  {32'hc26fa718, 32'h00000000} /* (13, 14, 16) {real, imag} */,
  {32'hc1a7668c, 32'hc1d67262} /* (13, 14, 15) {real, imag} */,
  {32'hc0c02acc, 32'hc0d97790} /* (13, 14, 14) {real, imag} */,
  {32'hc283eff7, 32'h41f7104c} /* (13, 14, 13) {real, imag} */,
  {32'h42c633ac, 32'h41b8b4ec} /* (13, 14, 12) {real, imag} */,
  {32'hc2aa5e58, 32'hc11a432c} /* (13, 14, 11) {real, imag} */,
  {32'hc26dfe05, 32'h4297bd1d} /* (13, 14, 10) {real, imag} */,
  {32'hc220d328, 32'hc1485a27} /* (13, 14, 9) {real, imag} */,
  {32'h4057b9a0, 32'h41c6fae8} /* (13, 14, 8) {real, imag} */,
  {32'hc2facc9e, 32'h42aacad4} /* (13, 14, 7) {real, imag} */,
  {32'h4034c520, 32'h433bb03f} /* (13, 14, 6) {real, imag} */,
  {32'h42a6d26c, 32'h42f14d76} /* (13, 14, 5) {real, imag} */,
  {32'hc314b843, 32'hc2807fd0} /* (13, 14, 4) {real, imag} */,
  {32'h413c3e48, 32'h41e4a0ea} /* (13, 14, 3) {real, imag} */,
  {32'h44839641, 32'h43457762} /* (13, 14, 2) {real, imag} */,
  {32'hc551ba7e, 32'hc3813898} /* (13, 14, 1) {real, imag} */,
  {32'hc50f0074, 32'h00000000} /* (13, 14, 0) {real, imag} */,
  {32'hc533aec8, 32'h4336a98c} /* (13, 13, 31) {real, imag} */,
  {32'h447c793e, 32'hc30f8d31} /* (13, 13, 30) {real, imag} */,
  {32'h42847450, 32'h4293e452} /* (13, 13, 29) {real, imag} */,
  {32'hc303b72c, 32'h4306f499} /* (13, 13, 28) {real, imag} */,
  {32'h42968b76, 32'hc2b9e43c} /* (13, 13, 27) {real, imag} */,
  {32'h41b77b91, 32'hc2cea07e} /* (13, 13, 26) {real, imag} */,
  {32'h41faaad5, 32'h3fcb99c8} /* (13, 13, 25) {real, imag} */,
  {32'hc2788a0b, 32'hc1eddf67} /* (13, 13, 24) {real, imag} */,
  {32'h4206295f, 32'h42948eb8} /* (13, 13, 23) {real, imag} */,
  {32'hc1dd8e53, 32'hc284092d} /* (13, 13, 22) {real, imag} */,
  {32'h423c3a04, 32'hc3026bf4} /* (13, 13, 21) {real, imag} */,
  {32'hc1c5e5fc, 32'h4145a940} /* (13, 13, 20) {real, imag} */,
  {32'hc1f5c558, 32'h41f21ac0} /* (13, 13, 19) {real, imag} */,
  {32'hc24355af, 32'h41a3dbe2} /* (13, 13, 18) {real, imag} */,
  {32'h41ec049a, 32'hc1ed5135} /* (13, 13, 17) {real, imag} */,
  {32'hc199b4f2, 32'h00000000} /* (13, 13, 16) {real, imag} */,
  {32'h41ec049a, 32'h41ed5135} /* (13, 13, 15) {real, imag} */,
  {32'hc24355af, 32'hc1a3dbe2} /* (13, 13, 14) {real, imag} */,
  {32'hc1f5c558, 32'hc1f21ac0} /* (13, 13, 13) {real, imag} */,
  {32'hc1c5e5fc, 32'hc145a940} /* (13, 13, 12) {real, imag} */,
  {32'h423c3a04, 32'h43026bf4} /* (13, 13, 11) {real, imag} */,
  {32'hc1dd8e53, 32'h4284092d} /* (13, 13, 10) {real, imag} */,
  {32'h4206295f, 32'hc2948eb8} /* (13, 13, 9) {real, imag} */,
  {32'hc2788a0b, 32'h41eddf67} /* (13, 13, 8) {real, imag} */,
  {32'h41faaad5, 32'hbfcb99c8} /* (13, 13, 7) {real, imag} */,
  {32'h41b77b91, 32'h42cea07e} /* (13, 13, 6) {real, imag} */,
  {32'h42968b76, 32'h42b9e43c} /* (13, 13, 5) {real, imag} */,
  {32'hc303b72c, 32'hc306f499} /* (13, 13, 4) {real, imag} */,
  {32'h42847450, 32'hc293e452} /* (13, 13, 3) {real, imag} */,
  {32'h447c793e, 32'h430f8d31} /* (13, 13, 2) {real, imag} */,
  {32'hc533aec8, 32'hc336a98c} /* (13, 13, 1) {real, imag} */,
  {32'hc4e0a9a2, 32'h00000000} /* (13, 13, 0) {real, imag} */,
  {32'hc5112cee, 32'h424229b0} /* (13, 12, 31) {real, imag} */,
  {32'h444aa16a, 32'h411a2190} /* (13, 12, 30) {real, imag} */,
  {32'h42fbe731, 32'h42212043} /* (13, 12, 29) {real, imag} */,
  {32'hc3281aae, 32'h438e8584} /* (13, 12, 28) {real, imag} */,
  {32'h437a9bd6, 32'hc2f5c150} /* (13, 12, 27) {real, imag} */,
  {32'h42e7dbfe, 32'hc2dd8428} /* (13, 12, 26) {real, imag} */,
  {32'hc19a5d58, 32'h41c4e8da} /* (13, 12, 25) {real, imag} */,
  {32'h42aca27a, 32'hc3660848} /* (13, 12, 24) {real, imag} */,
  {32'hc26d1090, 32'h42f9917f} /* (13, 12, 23) {real, imag} */,
  {32'hc1d88568, 32'hc13e289a} /* (13, 12, 22) {real, imag} */,
  {32'h41444d60, 32'h41c10fe6} /* (13, 12, 21) {real, imag} */,
  {32'h41af70f6, 32'h42bc5cf4} /* (13, 12, 20) {real, imag} */,
  {32'hc2617f84, 32'hc1f5aa52} /* (13, 12, 19) {real, imag} */,
  {32'hc24199c2, 32'hc15755de} /* (13, 12, 18) {real, imag} */,
  {32'h42804114, 32'hc248552f} /* (13, 12, 17) {real, imag} */,
  {32'h416c656a, 32'h00000000} /* (13, 12, 16) {real, imag} */,
  {32'h42804114, 32'h4248552f} /* (13, 12, 15) {real, imag} */,
  {32'hc24199c2, 32'h415755de} /* (13, 12, 14) {real, imag} */,
  {32'hc2617f84, 32'h41f5aa52} /* (13, 12, 13) {real, imag} */,
  {32'h41af70f6, 32'hc2bc5cf4} /* (13, 12, 12) {real, imag} */,
  {32'h41444d60, 32'hc1c10fe6} /* (13, 12, 11) {real, imag} */,
  {32'hc1d88568, 32'h413e289a} /* (13, 12, 10) {real, imag} */,
  {32'hc26d1090, 32'hc2f9917f} /* (13, 12, 9) {real, imag} */,
  {32'h42aca27a, 32'h43660848} /* (13, 12, 8) {real, imag} */,
  {32'hc19a5d58, 32'hc1c4e8da} /* (13, 12, 7) {real, imag} */,
  {32'h42e7dbfe, 32'h42dd8428} /* (13, 12, 6) {real, imag} */,
  {32'h437a9bd6, 32'h42f5c150} /* (13, 12, 5) {real, imag} */,
  {32'hc3281aae, 32'hc38e8584} /* (13, 12, 4) {real, imag} */,
  {32'h42fbe731, 32'hc2212043} /* (13, 12, 3) {real, imag} */,
  {32'h444aa16a, 32'hc11a2190} /* (13, 12, 2) {real, imag} */,
  {32'hc5112cee, 32'hc24229b0} /* (13, 12, 1) {real, imag} */,
  {32'hc48607fd, 32'h00000000} /* (13, 12, 0) {real, imag} */,
  {32'hc4a00a02, 32'hc352bcb4} /* (13, 11, 31) {real, imag} */,
  {32'h440e621e, 32'hc1dcac58} /* (13, 11, 30) {real, imag} */,
  {32'h42aead44, 32'h4293d19c} /* (13, 11, 29) {real, imag} */,
  {32'hc2cb7a57, 32'h43227f78} /* (13, 11, 28) {real, imag} */,
  {32'h4248e170, 32'hc31973ac} /* (13, 11, 27) {real, imag} */,
  {32'h425de284, 32'h423b5646} /* (13, 11, 26) {real, imag} */,
  {32'hc2ba5231, 32'hc309c449} /* (13, 11, 25) {real, imag} */,
  {32'h42973328, 32'h42217d5d} /* (13, 11, 24) {real, imag} */,
  {32'h41adf052, 32'h42d71394} /* (13, 11, 23) {real, imag} */,
  {32'hc2b0e89f, 32'h42ac127c} /* (13, 11, 22) {real, imag} */,
  {32'hc28e315e, 32'hc29097a4} /* (13, 11, 21) {real, imag} */,
  {32'h421c5ecb, 32'hc15ab03a} /* (13, 11, 20) {real, imag} */,
  {32'h4293a6dd, 32'hc2843cb8} /* (13, 11, 19) {real, imag} */,
  {32'h4204b3fa, 32'hc29be80a} /* (13, 11, 18) {real, imag} */,
  {32'hc23da60e, 32'h4171f660} /* (13, 11, 17) {real, imag} */,
  {32'hc2c2ac4b, 32'h00000000} /* (13, 11, 16) {real, imag} */,
  {32'hc23da60e, 32'hc171f660} /* (13, 11, 15) {real, imag} */,
  {32'h4204b3fa, 32'h429be80a} /* (13, 11, 14) {real, imag} */,
  {32'h4293a6dd, 32'h42843cb8} /* (13, 11, 13) {real, imag} */,
  {32'h421c5ecb, 32'h415ab03a} /* (13, 11, 12) {real, imag} */,
  {32'hc28e315e, 32'h429097a4} /* (13, 11, 11) {real, imag} */,
  {32'hc2b0e89f, 32'hc2ac127c} /* (13, 11, 10) {real, imag} */,
  {32'h41adf052, 32'hc2d71394} /* (13, 11, 9) {real, imag} */,
  {32'h42973328, 32'hc2217d5d} /* (13, 11, 8) {real, imag} */,
  {32'hc2ba5231, 32'h4309c449} /* (13, 11, 7) {real, imag} */,
  {32'h425de284, 32'hc23b5646} /* (13, 11, 6) {real, imag} */,
  {32'h4248e170, 32'h431973ac} /* (13, 11, 5) {real, imag} */,
  {32'hc2cb7a57, 32'hc3227f78} /* (13, 11, 4) {real, imag} */,
  {32'h42aead44, 32'hc293d19c} /* (13, 11, 3) {real, imag} */,
  {32'h440e621e, 32'h41dcac58} /* (13, 11, 2) {real, imag} */,
  {32'hc4a00a02, 32'h4352bcb4} /* (13, 11, 1) {real, imag} */,
  {32'hc350bd94, 32'h00000000} /* (13, 11, 0) {real, imag} */,
  {32'h43f2d436, 32'hc3e52bb4} /* (13, 10, 31) {real, imag} */,
  {32'h426c8090, 32'hc11300e0} /* (13, 10, 30) {real, imag} */,
  {32'hc2cd52ae, 32'hc1b92d46} /* (13, 10, 29) {real, imag} */,
  {32'h41ede728, 32'hc29d4182} /* (13, 10, 28) {real, imag} */,
  {32'hc2caa302, 32'hc2112e0c} /* (13, 10, 27) {real, imag} */,
  {32'hc2b0893a, 32'h426265f0} /* (13, 10, 26) {real, imag} */,
  {32'h420fd926, 32'hc2ba83a7} /* (13, 10, 25) {real, imag} */,
  {32'hc20c10a0, 32'h427f5894} /* (13, 10, 24) {real, imag} */,
  {32'h3f57bb00, 32'hc325ee10} /* (13, 10, 23) {real, imag} */,
  {32'h41a8f99f, 32'h418205ab} /* (13, 10, 22) {real, imag} */,
  {32'hc2be73b3, 32'hc27bef8f} /* (13, 10, 21) {real, imag} */,
  {32'hc2a900aa, 32'h423aee4d} /* (13, 10, 20) {real, imag} */,
  {32'h41beaef9, 32'hc18697b2} /* (13, 10, 19) {real, imag} */,
  {32'hc2dd5171, 32'h427fdcb4} /* (13, 10, 18) {real, imag} */,
  {32'h4240eaec, 32'h42a1b1df} /* (13, 10, 17) {real, imag} */,
  {32'hc110f4b6, 32'h00000000} /* (13, 10, 16) {real, imag} */,
  {32'h4240eaec, 32'hc2a1b1df} /* (13, 10, 15) {real, imag} */,
  {32'hc2dd5171, 32'hc27fdcb4} /* (13, 10, 14) {real, imag} */,
  {32'h41beaef9, 32'h418697b2} /* (13, 10, 13) {real, imag} */,
  {32'hc2a900aa, 32'hc23aee4d} /* (13, 10, 12) {real, imag} */,
  {32'hc2be73b3, 32'h427bef8f} /* (13, 10, 11) {real, imag} */,
  {32'h41a8f99f, 32'hc18205ab} /* (13, 10, 10) {real, imag} */,
  {32'h3f57bb00, 32'h4325ee10} /* (13, 10, 9) {real, imag} */,
  {32'hc20c10a0, 32'hc27f5894} /* (13, 10, 8) {real, imag} */,
  {32'h420fd926, 32'h42ba83a7} /* (13, 10, 7) {real, imag} */,
  {32'hc2b0893a, 32'hc26265f0} /* (13, 10, 6) {real, imag} */,
  {32'hc2caa302, 32'h42112e0c} /* (13, 10, 5) {real, imag} */,
  {32'h41ede728, 32'h429d4182} /* (13, 10, 4) {real, imag} */,
  {32'hc2cd52ae, 32'h41b92d46} /* (13, 10, 3) {real, imag} */,
  {32'h426c8090, 32'h411300e0} /* (13, 10, 2) {real, imag} */,
  {32'h43f2d436, 32'h43e52bb4} /* (13, 10, 1) {real, imag} */,
  {32'h4483f277, 32'h00000000} /* (13, 10, 0) {real, imag} */,
  {32'h44c99f1e, 32'hc42b5b13} /* (13, 9, 31) {real, imag} */,
  {32'hc4311026, 32'h438ca72c} /* (13, 9, 30) {real, imag} */,
  {32'hc2a50862, 32'h41aefd5c} /* (13, 9, 29) {real, imag} */,
  {32'h42164af2, 32'h41c561d8} /* (13, 9, 28) {real, imag} */,
  {32'hc2a9b058, 32'h4243fea8} /* (13, 9, 27) {real, imag} */,
  {32'h40d47ea8, 32'hc094a704} /* (13, 9, 26) {real, imag} */,
  {32'h429ae296, 32'h4250a77e} /* (13, 9, 25) {real, imag} */,
  {32'h42819444, 32'h41f2a8e8} /* (13, 9, 24) {real, imag} */,
  {32'h41013244, 32'h407f19b0} /* (13, 9, 23) {real, imag} */,
  {32'hc195868e, 32'hc2620c2b} /* (13, 9, 22) {real, imag} */,
  {32'hc2f772a8, 32'h42fc0f0e} /* (13, 9, 21) {real, imag} */,
  {32'h42148d92, 32'hc2c8cca0} /* (13, 9, 20) {real, imag} */,
  {32'h43103c51, 32'hc1d4a0bc} /* (13, 9, 19) {real, imag} */,
  {32'hc2aa03d1, 32'h429ed6db} /* (13, 9, 18) {real, imag} */,
  {32'h42bd44d0, 32'h421a07da} /* (13, 9, 17) {real, imag} */,
  {32'hc2c249b9, 32'h00000000} /* (13, 9, 16) {real, imag} */,
  {32'h42bd44d0, 32'hc21a07da} /* (13, 9, 15) {real, imag} */,
  {32'hc2aa03d1, 32'hc29ed6db} /* (13, 9, 14) {real, imag} */,
  {32'h43103c51, 32'h41d4a0bc} /* (13, 9, 13) {real, imag} */,
  {32'h42148d92, 32'h42c8cca0} /* (13, 9, 12) {real, imag} */,
  {32'hc2f772a8, 32'hc2fc0f0e} /* (13, 9, 11) {real, imag} */,
  {32'hc195868e, 32'h42620c2b} /* (13, 9, 10) {real, imag} */,
  {32'h41013244, 32'hc07f19b0} /* (13, 9, 9) {real, imag} */,
  {32'h42819444, 32'hc1f2a8e8} /* (13, 9, 8) {real, imag} */,
  {32'h429ae296, 32'hc250a77e} /* (13, 9, 7) {real, imag} */,
  {32'h40d47ea8, 32'h4094a704} /* (13, 9, 6) {real, imag} */,
  {32'hc2a9b058, 32'hc243fea8} /* (13, 9, 5) {real, imag} */,
  {32'h42164af2, 32'hc1c561d8} /* (13, 9, 4) {real, imag} */,
  {32'hc2a50862, 32'hc1aefd5c} /* (13, 9, 3) {real, imag} */,
  {32'hc4311026, 32'hc38ca72c} /* (13, 9, 2) {real, imag} */,
  {32'h44c99f1e, 32'h442b5b13} /* (13, 9, 1) {real, imag} */,
  {32'h44f6d6b0, 32'h00000000} /* (13, 9, 0) {real, imag} */,
  {32'h4509b4e7, 32'hc452f380} /* (13, 8, 31) {real, imag} */,
  {32'hc456ed5e, 32'h43e9d665} /* (13, 8, 30) {real, imag} */,
  {32'hc2b50594, 32'h4202408e} /* (13, 8, 29) {real, imag} */,
  {32'h43038ce6, 32'h417b9ee4} /* (13, 8, 28) {real, imag} */,
  {32'hc2a8c523, 32'h42af28d2} /* (13, 8, 27) {real, imag} */,
  {32'hc217ab99, 32'h42779ea8} /* (13, 8, 26) {real, imag} */,
  {32'h414293c4, 32'hc2c8a8c7} /* (13, 8, 25) {real, imag} */,
  {32'hc1916c78, 32'h4286b3c9} /* (13, 8, 24) {real, imag} */,
  {32'hc2a79dda, 32'hc2e77c3a} /* (13, 8, 23) {real, imag} */,
  {32'hc2bdcb37, 32'hc1b93d37} /* (13, 8, 22) {real, imag} */,
  {32'hc15dcd48, 32'h4269ecb0} /* (13, 8, 21) {real, imag} */,
  {32'hc1e9ab98, 32'hc2535447} /* (13, 8, 20) {real, imag} */,
  {32'h4208ec76, 32'hc18c137a} /* (13, 8, 19) {real, imag} */,
  {32'h4221b9e4, 32'hc05a9988} /* (13, 8, 18) {real, imag} */,
  {32'h41426c48, 32'h41d5430b} /* (13, 8, 17) {real, imag} */,
  {32'h41f13f36, 32'h00000000} /* (13, 8, 16) {real, imag} */,
  {32'h41426c48, 32'hc1d5430b} /* (13, 8, 15) {real, imag} */,
  {32'h4221b9e4, 32'h405a9988} /* (13, 8, 14) {real, imag} */,
  {32'h4208ec76, 32'h418c137a} /* (13, 8, 13) {real, imag} */,
  {32'hc1e9ab98, 32'h42535447} /* (13, 8, 12) {real, imag} */,
  {32'hc15dcd48, 32'hc269ecb0} /* (13, 8, 11) {real, imag} */,
  {32'hc2bdcb37, 32'h41b93d37} /* (13, 8, 10) {real, imag} */,
  {32'hc2a79dda, 32'h42e77c3a} /* (13, 8, 9) {real, imag} */,
  {32'hc1916c78, 32'hc286b3c9} /* (13, 8, 8) {real, imag} */,
  {32'h414293c4, 32'h42c8a8c7} /* (13, 8, 7) {real, imag} */,
  {32'hc217ab99, 32'hc2779ea8} /* (13, 8, 6) {real, imag} */,
  {32'hc2a8c523, 32'hc2af28d2} /* (13, 8, 5) {real, imag} */,
  {32'h43038ce6, 32'hc17b9ee4} /* (13, 8, 4) {real, imag} */,
  {32'hc2b50594, 32'hc202408e} /* (13, 8, 3) {real, imag} */,
  {32'hc456ed5e, 32'hc3e9d665} /* (13, 8, 2) {real, imag} */,
  {32'h4509b4e7, 32'h4452f380} /* (13, 8, 1) {real, imag} */,
  {32'h45216ccc, 32'h00000000} /* (13, 8, 0) {real, imag} */,
  {32'h452068e2, 32'hc492fb18} /* (13, 7, 31) {real, imag} */,
  {32'hc4672d8c, 32'h441fc6a2} /* (13, 7, 30) {real, imag} */,
  {32'hc31398e4, 32'h4313a6bc} /* (13, 7, 29) {real, imag} */,
  {32'h4356d473, 32'hc31acee6} /* (13, 7, 28) {real, imag} */,
  {32'hc346aa70, 32'h42e804d0} /* (13, 7, 27) {real, imag} */,
  {32'hc2269f70, 32'h43198cb0} /* (13, 7, 26) {real, imag} */,
  {32'h42963921, 32'hc2ee5ab5} /* (13, 7, 25) {real, imag} */,
  {32'hc2fad5db, 32'hc1117fcc} /* (13, 7, 24) {real, imag} */,
  {32'hc1210aac, 32'h40568f10} /* (13, 7, 23) {real, imag} */,
  {32'h42a08e80, 32'h40837908} /* (13, 7, 22) {real, imag} */,
  {32'hc2f8ba2e, 32'h43262ab2} /* (13, 7, 21) {real, imag} */,
  {32'hc15edd4a, 32'hc2753cd7} /* (13, 7, 20) {real, imag} */,
  {32'hc195a992, 32'hc29b1eb1} /* (13, 7, 19) {real, imag} */,
  {32'hc0790018, 32'h4200d682} /* (13, 7, 18) {real, imag} */,
  {32'hc0e8bbf0, 32'h42953000} /* (13, 7, 17) {real, imag} */,
  {32'h4211d12a, 32'h00000000} /* (13, 7, 16) {real, imag} */,
  {32'hc0e8bbf0, 32'hc2953000} /* (13, 7, 15) {real, imag} */,
  {32'hc0790018, 32'hc200d682} /* (13, 7, 14) {real, imag} */,
  {32'hc195a992, 32'h429b1eb1} /* (13, 7, 13) {real, imag} */,
  {32'hc15edd4a, 32'h42753cd7} /* (13, 7, 12) {real, imag} */,
  {32'hc2f8ba2e, 32'hc3262ab2} /* (13, 7, 11) {real, imag} */,
  {32'h42a08e80, 32'hc0837908} /* (13, 7, 10) {real, imag} */,
  {32'hc1210aac, 32'hc0568f10} /* (13, 7, 9) {real, imag} */,
  {32'hc2fad5db, 32'h41117fcc} /* (13, 7, 8) {real, imag} */,
  {32'h42963921, 32'h42ee5ab5} /* (13, 7, 7) {real, imag} */,
  {32'hc2269f70, 32'hc3198cb0} /* (13, 7, 6) {real, imag} */,
  {32'hc346aa70, 32'hc2e804d0} /* (13, 7, 5) {real, imag} */,
  {32'h4356d473, 32'h431acee6} /* (13, 7, 4) {real, imag} */,
  {32'hc31398e4, 32'hc313a6bc} /* (13, 7, 3) {real, imag} */,
  {32'hc4672d8c, 32'hc41fc6a2} /* (13, 7, 2) {real, imag} */,
  {32'h452068e2, 32'h4492fb18} /* (13, 7, 1) {real, imag} */,
  {32'h453d0a14, 32'h00000000} /* (13, 7, 0) {real, imag} */,
  {32'h4522b7fa, 32'hc4d1e92e} /* (13, 6, 31) {real, imag} */,
  {32'hc4442454, 32'h442d64c8} /* (13, 6, 30) {real, imag} */,
  {32'hc2e9a58a, 32'h42c5702a} /* (13, 6, 29) {real, imag} */,
  {32'h428a18d2, 32'hc2fe6a62} /* (13, 6, 28) {real, imag} */,
  {32'hc32c7636, 32'h43202db7} /* (13, 6, 27) {real, imag} */,
  {32'h42990362, 32'h41ee17dd} /* (13, 6, 26) {real, imag} */,
  {32'h41c614b5, 32'hc1ddffaa} /* (13, 6, 25) {real, imag} */,
  {32'hc1b6b30c, 32'h4108a008} /* (13, 6, 24) {real, imag} */,
  {32'h42ba350a, 32'hc1deb4c3} /* (13, 6, 23) {real, imag} */,
  {32'hc1660b2c, 32'hc262c020} /* (13, 6, 22) {real, imag} */,
  {32'hc2b36d8a, 32'h422ebc56} /* (13, 6, 21) {real, imag} */,
  {32'hc21797fc, 32'h428cd5dc} /* (13, 6, 20) {real, imag} */,
  {32'hc181bbd5, 32'hc201b1f8} /* (13, 6, 19) {real, imag} */,
  {32'h418adbed, 32'hc201e4a4} /* (13, 6, 18) {real, imag} */,
  {32'h41074ad8, 32'hc2929c61} /* (13, 6, 17) {real, imag} */,
  {32'h41dcf287, 32'h00000000} /* (13, 6, 16) {real, imag} */,
  {32'h41074ad8, 32'h42929c61} /* (13, 6, 15) {real, imag} */,
  {32'h418adbed, 32'h4201e4a4} /* (13, 6, 14) {real, imag} */,
  {32'hc181bbd5, 32'h4201b1f8} /* (13, 6, 13) {real, imag} */,
  {32'hc21797fc, 32'hc28cd5dc} /* (13, 6, 12) {real, imag} */,
  {32'hc2b36d8a, 32'hc22ebc56} /* (13, 6, 11) {real, imag} */,
  {32'hc1660b2c, 32'h4262c020} /* (13, 6, 10) {real, imag} */,
  {32'h42ba350a, 32'h41deb4c3} /* (13, 6, 9) {real, imag} */,
  {32'hc1b6b30c, 32'hc108a008} /* (13, 6, 8) {real, imag} */,
  {32'h41c614b5, 32'h41ddffaa} /* (13, 6, 7) {real, imag} */,
  {32'h42990362, 32'hc1ee17dd} /* (13, 6, 6) {real, imag} */,
  {32'hc32c7636, 32'hc3202db7} /* (13, 6, 5) {real, imag} */,
  {32'h428a18d2, 32'h42fe6a62} /* (13, 6, 4) {real, imag} */,
  {32'hc2e9a58a, 32'hc2c5702a} /* (13, 6, 3) {real, imag} */,
  {32'hc4442454, 32'hc42d64c8} /* (13, 6, 2) {real, imag} */,
  {32'h4522b7fa, 32'h44d1e92e} /* (13, 6, 1) {real, imag} */,
  {32'h45571d72, 32'h00000000} /* (13, 6, 0) {real, imag} */,
  {32'h451b783c, 32'hc513e397} /* (13, 5, 31) {real, imag} */,
  {32'hc33a40d8, 32'h445234ff} /* (13, 5, 30) {real, imag} */,
  {32'hc30bb87a, 32'h4253be3a} /* (13, 5, 29) {real, imag} */,
  {32'hc305fe5d, 32'h428f0591} /* (13, 5, 28) {real, imag} */,
  {32'hc34641ab, 32'hc18c2a8c} /* (13, 5, 27) {real, imag} */,
  {32'h4312ee3b, 32'h4122eb4f} /* (13, 5, 26) {real, imag} */,
  {32'hc205b59c, 32'hc2cf5146} /* (13, 5, 25) {real, imag} */,
  {32'hc10ae21c, 32'h4315cd25} /* (13, 5, 24) {real, imag} */,
  {32'hc2827a76, 32'hc2416b2a} /* (13, 5, 23) {real, imag} */,
  {32'hc1f46296, 32'h41cdb22a} /* (13, 5, 22) {real, imag} */,
  {32'h40a7f000, 32'h41bcc153} /* (13, 5, 21) {real, imag} */,
  {32'h425ca67c, 32'h41e70e5c} /* (13, 5, 20) {real, imag} */,
  {32'h420bc30c, 32'hc0a8b360} /* (13, 5, 19) {real, imag} */,
  {32'hc24464f9, 32'h4172f81d} /* (13, 5, 18) {real, imag} */,
  {32'h41baf0db, 32'hc21106b6} /* (13, 5, 17) {real, imag} */,
  {32'hc30e8202, 32'h00000000} /* (13, 5, 16) {real, imag} */,
  {32'h41baf0db, 32'h421106b6} /* (13, 5, 15) {real, imag} */,
  {32'hc24464f9, 32'hc172f81d} /* (13, 5, 14) {real, imag} */,
  {32'h420bc30c, 32'h40a8b360} /* (13, 5, 13) {real, imag} */,
  {32'h425ca67c, 32'hc1e70e5c} /* (13, 5, 12) {real, imag} */,
  {32'h40a7f000, 32'hc1bcc153} /* (13, 5, 11) {real, imag} */,
  {32'hc1f46296, 32'hc1cdb22a} /* (13, 5, 10) {real, imag} */,
  {32'hc2827a76, 32'h42416b2a} /* (13, 5, 9) {real, imag} */,
  {32'hc10ae21c, 32'hc315cd25} /* (13, 5, 8) {real, imag} */,
  {32'hc205b59c, 32'h42cf5146} /* (13, 5, 7) {real, imag} */,
  {32'h4312ee3b, 32'hc122eb4f} /* (13, 5, 6) {real, imag} */,
  {32'hc34641ab, 32'h418c2a8c} /* (13, 5, 5) {real, imag} */,
  {32'hc305fe5d, 32'hc28f0591} /* (13, 5, 4) {real, imag} */,
  {32'hc30bb87a, 32'hc253be3a} /* (13, 5, 3) {real, imag} */,
  {32'hc33a40d8, 32'hc45234ff} /* (13, 5, 2) {real, imag} */,
  {32'h451b783c, 32'h4513e397} /* (13, 5, 1) {real, imag} */,
  {32'h456c3f1f, 32'h00000000} /* (13, 5, 0) {real, imag} */,
  {32'h450e485a, 32'hc53b300e} /* (13, 4, 31) {real, imag} */,
  {32'h42fe2590, 32'h448a3ed4} /* (13, 4, 30) {real, imag} */,
  {32'hc26820a0, 32'h42ca6ca4} /* (13, 4, 29) {real, imag} */,
  {32'hc32aed44, 32'h42669064} /* (13, 4, 28) {real, imag} */,
  {32'hc38067aa, 32'hc2a390a6} /* (13, 4, 27) {real, imag} */,
  {32'h42d37ca1, 32'h42b7cc38} /* (13, 4, 26) {real, imag} */,
  {32'hc2b8b890, 32'hc2ccd902} /* (13, 4, 25) {real, imag} */,
  {32'h41f5cec9, 32'h42af3f3b} /* (13, 4, 24) {real, imag} */,
  {32'hc1fd8574, 32'h419537b5} /* (13, 4, 23) {real, imag} */,
  {32'hc1b7a222, 32'h418d68c4} /* (13, 4, 22) {real, imag} */,
  {32'hc1d68a2f, 32'hc226e0ad} /* (13, 4, 21) {real, imag} */,
  {32'h4289e5d8, 32'hc246b407} /* (13, 4, 20) {real, imag} */,
  {32'hc2456a5f, 32'h41e335c0} /* (13, 4, 19) {real, imag} */,
  {32'h4260f924, 32'hc264e228} /* (13, 4, 18) {real, imag} */,
  {32'hc19c0b65, 32'h41f79544} /* (13, 4, 17) {real, imag} */,
  {32'hc28b682f, 32'h00000000} /* (13, 4, 16) {real, imag} */,
  {32'hc19c0b65, 32'hc1f79544} /* (13, 4, 15) {real, imag} */,
  {32'h4260f924, 32'h4264e228} /* (13, 4, 14) {real, imag} */,
  {32'hc2456a5f, 32'hc1e335c0} /* (13, 4, 13) {real, imag} */,
  {32'h4289e5d8, 32'h4246b407} /* (13, 4, 12) {real, imag} */,
  {32'hc1d68a2f, 32'h4226e0ad} /* (13, 4, 11) {real, imag} */,
  {32'hc1b7a222, 32'hc18d68c4} /* (13, 4, 10) {real, imag} */,
  {32'hc1fd8574, 32'hc19537b5} /* (13, 4, 9) {real, imag} */,
  {32'h41f5cec9, 32'hc2af3f3b} /* (13, 4, 8) {real, imag} */,
  {32'hc2b8b890, 32'h42ccd902} /* (13, 4, 7) {real, imag} */,
  {32'h42d37ca1, 32'hc2b7cc38} /* (13, 4, 6) {real, imag} */,
  {32'hc38067aa, 32'h42a390a6} /* (13, 4, 5) {real, imag} */,
  {32'hc32aed44, 32'hc2669064} /* (13, 4, 4) {real, imag} */,
  {32'hc26820a0, 32'hc2ca6ca4} /* (13, 4, 3) {real, imag} */,
  {32'h42fe2590, 32'hc48a3ed4} /* (13, 4, 2) {real, imag} */,
  {32'h450e485a, 32'h453b300e} /* (13, 4, 1) {real, imag} */,
  {32'h45822e7f, 32'h00000000} /* (13, 4, 0) {real, imag} */,
  {32'h4516776d, 32'hc54611c2} /* (13, 3, 31) {real, imag} */,
  {32'h42afdb30, 32'h44866c82} /* (13, 3, 30) {real, imag} */,
  {32'hc376639f, 32'h431d58f3} /* (13, 3, 29) {real, imag} */,
  {32'hc27f020f, 32'h42a90fd7} /* (13, 3, 28) {real, imag} */,
  {32'hc31b40df, 32'hc29be44e} /* (13, 3, 27) {real, imag} */,
  {32'h419a7710, 32'h416f3130} /* (13, 3, 26) {real, imag} */,
  {32'h4280adb9, 32'hc2ba4074} /* (13, 3, 25) {real, imag} */,
  {32'h42eab7b0, 32'h41adc308} /* (13, 3, 24) {real, imag} */,
  {32'h4282bb4b, 32'hc2b0459e} /* (13, 3, 23) {real, imag} */,
  {32'hc23f4619, 32'h4219e218} /* (13, 3, 22) {real, imag} */,
  {32'hc215ca34, 32'h430327a1} /* (13, 3, 21) {real, imag} */,
  {32'hc21ba82c, 32'hc205c600} /* (13, 3, 20) {real, imag} */,
  {32'h429a7e5a, 32'hc2292563} /* (13, 3, 19) {real, imag} */,
  {32'hc2a41618, 32'h42ae9c3a} /* (13, 3, 18) {real, imag} */,
  {32'h41937db2, 32'hc23979d6} /* (13, 3, 17) {real, imag} */,
  {32'h431e4310, 32'h00000000} /* (13, 3, 16) {real, imag} */,
  {32'h41937db2, 32'h423979d6} /* (13, 3, 15) {real, imag} */,
  {32'hc2a41618, 32'hc2ae9c3a} /* (13, 3, 14) {real, imag} */,
  {32'h429a7e5a, 32'h42292563} /* (13, 3, 13) {real, imag} */,
  {32'hc21ba82c, 32'h4205c600} /* (13, 3, 12) {real, imag} */,
  {32'hc215ca34, 32'hc30327a1} /* (13, 3, 11) {real, imag} */,
  {32'hc23f4619, 32'hc219e218} /* (13, 3, 10) {real, imag} */,
  {32'h4282bb4b, 32'h42b0459e} /* (13, 3, 9) {real, imag} */,
  {32'h42eab7b0, 32'hc1adc308} /* (13, 3, 8) {real, imag} */,
  {32'h4280adb9, 32'h42ba4074} /* (13, 3, 7) {real, imag} */,
  {32'h419a7710, 32'hc16f3130} /* (13, 3, 6) {real, imag} */,
  {32'hc31b40df, 32'h429be44e} /* (13, 3, 5) {real, imag} */,
  {32'hc27f020f, 32'hc2a90fd7} /* (13, 3, 4) {real, imag} */,
  {32'hc376639f, 32'hc31d58f3} /* (13, 3, 3) {real, imag} */,
  {32'h42afdb30, 32'hc4866c82} /* (13, 3, 2) {real, imag} */,
  {32'h4516776d, 32'h454611c2} /* (13, 3, 1) {real, imag} */,
  {32'h4581e5f3, 32'h00000000} /* (13, 3, 0) {real, imag} */,
  {32'h451b704e, 32'hc543605f} /* (13, 2, 31) {real, imag} */,
  {32'h42d68090, 32'h44582af8} /* (13, 2, 30) {real, imag} */,
  {32'hc38de468, 32'h43130b33} /* (13, 2, 29) {real, imag} */,
  {32'hc3375759, 32'h4356c2d2} /* (13, 2, 28) {real, imag} */,
  {32'hc32ae879, 32'hc3148a6a} /* (13, 2, 27) {real, imag} */,
  {32'h41e991c8, 32'h41503c58} /* (13, 2, 26) {real, imag} */,
  {32'hc1c8800e, 32'h426ac5e0} /* (13, 2, 25) {real, imag} */,
  {32'h42d9d028, 32'h42c3ef1a} /* (13, 2, 24) {real, imag} */,
  {32'hc2e6fa0e, 32'h428c9116} /* (13, 2, 23) {real, imag} */,
  {32'hc0d5b340, 32'hc10e9d28} /* (13, 2, 22) {real, imag} */,
  {32'hc25c77ce, 32'h4234c343} /* (13, 2, 21) {real, imag} */,
  {32'h42d5fd44, 32'hc311b75d} /* (13, 2, 20) {real, imag} */,
  {32'hc2170556, 32'hc2d9611b} /* (13, 2, 19) {real, imag} */,
  {32'hc23a7f2c, 32'hc1f2a282} /* (13, 2, 18) {real, imag} */,
  {32'h427c80fc, 32'h423a83d0} /* (13, 2, 17) {real, imag} */,
  {32'h425a0fde, 32'h00000000} /* (13, 2, 16) {real, imag} */,
  {32'h427c80fc, 32'hc23a83d0} /* (13, 2, 15) {real, imag} */,
  {32'hc23a7f2c, 32'h41f2a282} /* (13, 2, 14) {real, imag} */,
  {32'hc2170556, 32'h42d9611b} /* (13, 2, 13) {real, imag} */,
  {32'h42d5fd44, 32'h4311b75d} /* (13, 2, 12) {real, imag} */,
  {32'hc25c77ce, 32'hc234c343} /* (13, 2, 11) {real, imag} */,
  {32'hc0d5b340, 32'h410e9d28} /* (13, 2, 10) {real, imag} */,
  {32'hc2e6fa0e, 32'hc28c9116} /* (13, 2, 9) {real, imag} */,
  {32'h42d9d028, 32'hc2c3ef1a} /* (13, 2, 8) {real, imag} */,
  {32'hc1c8800e, 32'hc26ac5e0} /* (13, 2, 7) {real, imag} */,
  {32'h41e991c8, 32'hc1503c58} /* (13, 2, 6) {real, imag} */,
  {32'hc32ae879, 32'h43148a6a} /* (13, 2, 5) {real, imag} */,
  {32'hc3375759, 32'hc356c2d2} /* (13, 2, 4) {real, imag} */,
  {32'hc38de468, 32'hc3130b33} /* (13, 2, 3) {real, imag} */,
  {32'h42d68090, 32'hc4582af8} /* (13, 2, 2) {real, imag} */,
  {32'h451b704e, 32'h4543605f} /* (13, 2, 1) {real, imag} */,
  {32'h45851f8a, 32'h00000000} /* (13, 2, 0) {real, imag} */,
  {32'h45169a59, 32'hc5339fd1} /* (13, 1, 31) {real, imag} */,
  {32'h430fb7b0, 32'h444647b0} /* (13, 1, 30) {real, imag} */,
  {32'hc312fb81, 32'h42b25605} /* (13, 1, 29) {real, imag} */,
  {32'hc2eab47b, 32'h4357b9e9} /* (13, 1, 28) {real, imag} */,
  {32'hc35459fc, 32'hc20b68b4} /* (13, 1, 27) {real, imag} */,
  {32'h42681bd0, 32'hc1c151a8} /* (13, 1, 26) {real, imag} */,
  {32'h4205fae5, 32'h423f6334} /* (13, 1, 25) {real, imag} */,
  {32'h42d739e4, 32'h42533740} /* (13, 1, 24) {real, imag} */,
  {32'hc305df20, 32'h42eb8e86} /* (13, 1, 23) {real, imag} */,
  {32'hc26fc7c0, 32'h42d702f6} /* (13, 1, 22) {real, imag} */,
  {32'hc1b801d9, 32'hc316d1bb} /* (13, 1, 21) {real, imag} */,
  {32'h422ca888, 32'hc241e521} /* (13, 1, 20) {real, imag} */,
  {32'h41c4d943, 32'hc114f838} /* (13, 1, 19) {real, imag} */,
  {32'h429b4c78, 32'h42064dea} /* (13, 1, 18) {real, imag} */,
  {32'hc2656904, 32'h414e2ad2} /* (13, 1, 17) {real, imag} */,
  {32'hc2a61462, 32'h00000000} /* (13, 1, 16) {real, imag} */,
  {32'hc2656904, 32'hc14e2ad2} /* (13, 1, 15) {real, imag} */,
  {32'h429b4c78, 32'hc2064dea} /* (13, 1, 14) {real, imag} */,
  {32'h41c4d943, 32'h4114f838} /* (13, 1, 13) {real, imag} */,
  {32'h422ca888, 32'h4241e521} /* (13, 1, 12) {real, imag} */,
  {32'hc1b801d9, 32'h4316d1bb} /* (13, 1, 11) {real, imag} */,
  {32'hc26fc7c0, 32'hc2d702f6} /* (13, 1, 10) {real, imag} */,
  {32'hc305df20, 32'hc2eb8e86} /* (13, 1, 9) {real, imag} */,
  {32'h42d739e4, 32'hc2533740} /* (13, 1, 8) {real, imag} */,
  {32'h4205fae5, 32'hc23f6334} /* (13, 1, 7) {real, imag} */,
  {32'h42681bd0, 32'h41c151a8} /* (13, 1, 6) {real, imag} */,
  {32'hc35459fc, 32'h420b68b4} /* (13, 1, 5) {real, imag} */,
  {32'hc2eab47b, 32'hc357b9e9} /* (13, 1, 4) {real, imag} */,
  {32'hc312fb81, 32'hc2b25605} /* (13, 1, 3) {real, imag} */,
  {32'h430fb7b0, 32'hc44647b0} /* (13, 1, 2) {real, imag} */,
  {32'h45169a59, 32'h45339fd1} /* (13, 1, 1) {real, imag} */,
  {32'h45789eee, 32'h00000000} /* (13, 1, 0) {real, imag} */,
  {32'h451b2866, 32'hc514bc3c} /* (13, 0, 31) {real, imag} */,
  {32'hc3146fa4, 32'h44225e6a} /* (13, 0, 30) {real, imag} */,
  {32'hc28c6e1f, 32'h4176ed4c} /* (13, 0, 29) {real, imag} */,
  {32'hc27a4123, 32'h433f5a24} /* (13, 0, 28) {real, imag} */,
  {32'hc11f5f00, 32'h4118b4c4} /* (13, 0, 27) {real, imag} */,
  {32'hc19e7989, 32'h41c36d7f} /* (13, 0, 26) {real, imag} */,
  {32'h4299b581, 32'hc2c60eda} /* (13, 0, 25) {real, imag} */,
  {32'h42c33b48, 32'h416f7e6c} /* (13, 0, 24) {real, imag} */,
  {32'h416bfabc, 32'hc1861b3c} /* (13, 0, 23) {real, imag} */,
  {32'hc2298a9b, 32'h429081a4} /* (13, 0, 22) {real, imag} */,
  {32'h42ddf547, 32'hc203b44a} /* (13, 0, 21) {real, imag} */,
  {32'hc11ea800, 32'h4243ecf4} /* (13, 0, 20) {real, imag} */,
  {32'h4219aa53, 32'h4097ca2c} /* (13, 0, 19) {real, imag} */,
  {32'hc0d90132, 32'h41e9a982} /* (13, 0, 18) {real, imag} */,
  {32'h41b0b243, 32'h423f83c4} /* (13, 0, 17) {real, imag} */,
  {32'hc1fb8fa0, 32'h00000000} /* (13, 0, 16) {real, imag} */,
  {32'h41b0b243, 32'hc23f83c4} /* (13, 0, 15) {real, imag} */,
  {32'hc0d90132, 32'hc1e9a982} /* (13, 0, 14) {real, imag} */,
  {32'h4219aa53, 32'hc097ca2c} /* (13, 0, 13) {real, imag} */,
  {32'hc11ea800, 32'hc243ecf4} /* (13, 0, 12) {real, imag} */,
  {32'h42ddf547, 32'h4203b44a} /* (13, 0, 11) {real, imag} */,
  {32'hc2298a9b, 32'hc29081a4} /* (13, 0, 10) {real, imag} */,
  {32'h416bfabc, 32'h41861b3c} /* (13, 0, 9) {real, imag} */,
  {32'h42c33b48, 32'hc16f7e6c} /* (13, 0, 8) {real, imag} */,
  {32'h4299b581, 32'h42c60eda} /* (13, 0, 7) {real, imag} */,
  {32'hc19e7989, 32'hc1c36d7f} /* (13, 0, 6) {real, imag} */,
  {32'hc11f5f00, 32'hc118b4c4} /* (13, 0, 5) {real, imag} */,
  {32'hc27a4123, 32'hc33f5a24} /* (13, 0, 4) {real, imag} */,
  {32'hc28c6e1f, 32'hc176ed4c} /* (13, 0, 3) {real, imag} */,
  {32'hc3146fa4, 32'hc4225e6a} /* (13, 0, 2) {real, imag} */,
  {32'h451b2866, 32'h4514bc3c} /* (13, 0, 1) {real, imag} */,
  {32'h456f85db, 32'h00000000} /* (13, 0, 0) {real, imag} */,
  {32'h4562dca8, 32'hc4fe1114} /* (12, 31, 31) {real, imag} */,
  {32'hc43e1f30, 32'h4405257c} /* (12, 31, 30) {real, imag} */,
  {32'hc2e214d3, 32'h424782a0} /* (12, 31, 29) {real, imag} */,
  {32'h428011f0, 32'h42b31132} /* (12, 31, 28) {real, imag} */,
  {32'hc324e98e, 32'hc1363688} /* (12, 31, 27) {real, imag} */,
  {32'h426fd8a4, 32'hc0b4e7a6} /* (12, 31, 26) {real, imag} */,
  {32'hc1c0f072, 32'hc1e0f5d0} /* (12, 31, 25) {real, imag} */,
  {32'hc2d6702b, 32'h419b1306} /* (12, 31, 24) {real, imag} */,
  {32'hc25098ac, 32'hc14d36a4} /* (12, 31, 23) {real, imag} */,
  {32'h4192b884, 32'hc220775d} /* (12, 31, 22) {real, imag} */,
  {32'h419083be, 32'hc0063130} /* (12, 31, 21) {real, imag} */,
  {32'hc2611bd5, 32'hc2160a7a} /* (12, 31, 20) {real, imag} */,
  {32'hc11bf298, 32'hc23fb5d2} /* (12, 31, 19) {real, imag} */,
  {32'hc1ca0d17, 32'hc1b12e2b} /* (12, 31, 18) {real, imag} */,
  {32'h419fe09c, 32'h413887e5} /* (12, 31, 17) {real, imag} */,
  {32'h42960a7c, 32'h00000000} /* (12, 31, 16) {real, imag} */,
  {32'h419fe09c, 32'hc13887e5} /* (12, 31, 15) {real, imag} */,
  {32'hc1ca0d17, 32'h41b12e2b} /* (12, 31, 14) {real, imag} */,
  {32'hc11bf298, 32'h423fb5d2} /* (12, 31, 13) {real, imag} */,
  {32'hc2611bd5, 32'h42160a7a} /* (12, 31, 12) {real, imag} */,
  {32'h419083be, 32'h40063130} /* (12, 31, 11) {real, imag} */,
  {32'h4192b884, 32'h4220775d} /* (12, 31, 10) {real, imag} */,
  {32'hc25098ac, 32'h414d36a4} /* (12, 31, 9) {real, imag} */,
  {32'hc2d6702b, 32'hc19b1306} /* (12, 31, 8) {real, imag} */,
  {32'hc1c0f072, 32'h41e0f5d0} /* (12, 31, 7) {real, imag} */,
  {32'h426fd8a4, 32'h40b4e7a6} /* (12, 31, 6) {real, imag} */,
  {32'hc324e98e, 32'h41363688} /* (12, 31, 5) {real, imag} */,
  {32'h428011f0, 32'hc2b31132} /* (12, 31, 4) {real, imag} */,
  {32'hc2e214d3, 32'hc24782a0} /* (12, 31, 3) {real, imag} */,
  {32'hc43e1f30, 32'hc405257c} /* (12, 31, 2) {real, imag} */,
  {32'h4562dca8, 32'h44fe1114} /* (12, 31, 1) {real, imag} */,
  {32'h459754de, 32'h00000000} /* (12, 31, 0) {real, imag} */,
  {32'h45802c75, 32'hc4bb559a} /* (12, 30, 31) {real, imag} */,
  {32'hc49b914c, 32'h43fd5d01} /* (12, 30, 30) {real, imag} */,
  {32'h41f935f8, 32'h42ba8350} /* (12, 30, 29) {real, imag} */,
  {32'h429a323a, 32'hc25fb1a2} /* (12, 30, 28) {real, imag} */,
  {32'hc39594e0, 32'hc16f8608} /* (12, 30, 27) {real, imag} */,
  {32'h4220048d, 32'hc26959ca} /* (12, 30, 26) {real, imag} */,
  {32'h415bc9b8, 32'hc2cb1dc8} /* (12, 30, 25) {real, imag} */,
  {32'hc300eef4, 32'h412bfd04} /* (12, 30, 24) {real, imag} */,
  {32'hc23c2130, 32'hc1fdd50d} /* (12, 30, 23) {real, imag} */,
  {32'hc09bf254, 32'h4232701e} /* (12, 30, 22) {real, imag} */,
  {32'hc2ade723, 32'h40d48e4e} /* (12, 30, 21) {real, imag} */,
  {32'h3f2faf80, 32'h41ceaf39} /* (12, 30, 20) {real, imag} */,
  {32'h4285c932, 32'h41e6eb7c} /* (12, 30, 19) {real, imag} */,
  {32'h41211920, 32'hc23541d0} /* (12, 30, 18) {real, imag} */,
  {32'h4114ccfc, 32'h415ac87e} /* (12, 30, 17) {real, imag} */,
  {32'h42bdb6ce, 32'h00000000} /* (12, 30, 16) {real, imag} */,
  {32'h4114ccfc, 32'hc15ac87e} /* (12, 30, 15) {real, imag} */,
  {32'h41211920, 32'h423541d0} /* (12, 30, 14) {real, imag} */,
  {32'h4285c932, 32'hc1e6eb7c} /* (12, 30, 13) {real, imag} */,
  {32'h3f2faf80, 32'hc1ceaf39} /* (12, 30, 12) {real, imag} */,
  {32'hc2ade723, 32'hc0d48e4e} /* (12, 30, 11) {real, imag} */,
  {32'hc09bf254, 32'hc232701e} /* (12, 30, 10) {real, imag} */,
  {32'hc23c2130, 32'h41fdd50d} /* (12, 30, 9) {real, imag} */,
  {32'hc300eef4, 32'hc12bfd04} /* (12, 30, 8) {real, imag} */,
  {32'h415bc9b8, 32'h42cb1dc8} /* (12, 30, 7) {real, imag} */,
  {32'h4220048d, 32'h426959ca} /* (12, 30, 6) {real, imag} */,
  {32'hc39594e0, 32'h416f8608} /* (12, 30, 5) {real, imag} */,
  {32'h429a323a, 32'h425fb1a2} /* (12, 30, 4) {real, imag} */,
  {32'h41f935f8, 32'hc2ba8350} /* (12, 30, 3) {real, imag} */,
  {32'hc49b914c, 32'hc3fd5d01} /* (12, 30, 2) {real, imag} */,
  {32'h45802c75, 32'h44bb559a} /* (12, 30, 1) {real, imag} */,
  {32'h45a10627, 32'h00000000} /* (12, 30, 0) {real, imag} */,
  {32'h458d1089, 32'hc49f0e13} /* (12, 29, 31) {real, imag} */,
  {32'hc4bca606, 32'h43fa2828} /* (12, 29, 30) {real, imag} */,
  {32'h418a14a0, 32'h42b57ea2} /* (12, 29, 29) {real, imag} */,
  {32'h4303e162, 32'hc3449ba3} /* (12, 29, 28) {real, imag} */,
  {32'hc3687f36, 32'hc1f8ad50} /* (12, 29, 27) {real, imag} */,
  {32'h41dafbb6, 32'h4252ddba} /* (12, 29, 26) {real, imag} */,
  {32'hc2a166e6, 32'hc2377c3d} /* (12, 29, 25) {real, imag} */,
  {32'hc2ef8d02, 32'hc1cd0368} /* (12, 29, 24) {real, imag} */,
  {32'h40c530c2, 32'h40f92e30} /* (12, 29, 23) {real, imag} */,
  {32'hc1eeac34, 32'hc0865d80} /* (12, 29, 22) {real, imag} */,
  {32'h42770cce, 32'h41e27409} /* (12, 29, 21) {real, imag} */,
  {32'hc29be1e4, 32'h42c50a13} /* (12, 29, 20) {real, imag} */,
  {32'h427ac29f, 32'h42b81470} /* (12, 29, 19) {real, imag} */,
  {32'h4212da61, 32'h42af1ba8} /* (12, 29, 18) {real, imag} */,
  {32'hc121fdea, 32'h4064f560} /* (12, 29, 17) {real, imag} */,
  {32'hc25abac2, 32'h00000000} /* (12, 29, 16) {real, imag} */,
  {32'hc121fdea, 32'hc064f560} /* (12, 29, 15) {real, imag} */,
  {32'h4212da61, 32'hc2af1ba8} /* (12, 29, 14) {real, imag} */,
  {32'h427ac29f, 32'hc2b81470} /* (12, 29, 13) {real, imag} */,
  {32'hc29be1e4, 32'hc2c50a13} /* (12, 29, 12) {real, imag} */,
  {32'h42770cce, 32'hc1e27409} /* (12, 29, 11) {real, imag} */,
  {32'hc1eeac34, 32'h40865d80} /* (12, 29, 10) {real, imag} */,
  {32'h40c530c2, 32'hc0f92e30} /* (12, 29, 9) {real, imag} */,
  {32'hc2ef8d02, 32'h41cd0368} /* (12, 29, 8) {real, imag} */,
  {32'hc2a166e6, 32'h42377c3d} /* (12, 29, 7) {real, imag} */,
  {32'h41dafbb6, 32'hc252ddba} /* (12, 29, 6) {real, imag} */,
  {32'hc3687f36, 32'h41f8ad50} /* (12, 29, 5) {real, imag} */,
  {32'h4303e162, 32'h43449ba3} /* (12, 29, 4) {real, imag} */,
  {32'h418a14a0, 32'hc2b57ea2} /* (12, 29, 3) {real, imag} */,
  {32'hc4bca606, 32'hc3fa2828} /* (12, 29, 2) {real, imag} */,
  {32'h458d1089, 32'h449f0e13} /* (12, 29, 1) {real, imag} */,
  {32'h45a09f1d, 32'h00000000} /* (12, 29, 0) {real, imag} */,
  {32'h45977443, 32'hc48aead2} /* (12, 28, 31) {real, imag} */,
  {32'hc4ca5662, 32'h4392cd8a} /* (12, 28, 30) {real, imag} */,
  {32'hc2590de3, 32'h428696a6} /* (12, 28, 29) {real, imag} */,
  {32'h4307d336, 32'hc36c589d} /* (12, 28, 28) {real, imag} */,
  {32'hc351146d, 32'h420c5081} /* (12, 28, 27) {real, imag} */,
  {32'hc12562bd, 32'hc1f7980f} /* (12, 28, 26) {real, imag} */,
  {32'hc0644350, 32'h4270df96} /* (12, 28, 25) {real, imag} */,
  {32'hc2ffd0cd, 32'h41e1b714} /* (12, 28, 24) {real, imag} */,
  {32'hc06959d0, 32'h42ff780c} /* (12, 28, 23) {real, imag} */,
  {32'hc1208d60, 32'h430ff931} /* (12, 28, 22) {real, imag} */,
  {32'h428726db, 32'h42265d25} /* (12, 28, 21) {real, imag} */,
  {32'hc21255b9, 32'h40d1ac1c} /* (12, 28, 20) {real, imag} */,
  {32'hc2fc743a, 32'hc1fa9714} /* (12, 28, 19) {real, imag} */,
  {32'h4241ec22, 32'hc1aad4ec} /* (12, 28, 18) {real, imag} */,
  {32'h42a261d4, 32'hc29af4cc} /* (12, 28, 17) {real, imag} */,
  {32'h41e20aa2, 32'h00000000} /* (12, 28, 16) {real, imag} */,
  {32'h42a261d4, 32'h429af4cc} /* (12, 28, 15) {real, imag} */,
  {32'h4241ec22, 32'h41aad4ec} /* (12, 28, 14) {real, imag} */,
  {32'hc2fc743a, 32'h41fa9714} /* (12, 28, 13) {real, imag} */,
  {32'hc21255b9, 32'hc0d1ac1c} /* (12, 28, 12) {real, imag} */,
  {32'h428726db, 32'hc2265d25} /* (12, 28, 11) {real, imag} */,
  {32'hc1208d60, 32'hc30ff931} /* (12, 28, 10) {real, imag} */,
  {32'hc06959d0, 32'hc2ff780c} /* (12, 28, 9) {real, imag} */,
  {32'hc2ffd0cd, 32'hc1e1b714} /* (12, 28, 8) {real, imag} */,
  {32'hc0644350, 32'hc270df96} /* (12, 28, 7) {real, imag} */,
  {32'hc12562bd, 32'h41f7980f} /* (12, 28, 6) {real, imag} */,
  {32'hc351146d, 32'hc20c5081} /* (12, 28, 5) {real, imag} */,
  {32'h4307d336, 32'h436c589d} /* (12, 28, 4) {real, imag} */,
  {32'hc2590de3, 32'hc28696a6} /* (12, 28, 3) {real, imag} */,
  {32'hc4ca5662, 32'hc392cd8a} /* (12, 28, 2) {real, imag} */,
  {32'h45977443, 32'h448aead2} /* (12, 28, 1) {real, imag} */,
  {32'h459baf19, 32'h00000000} /* (12, 28, 0) {real, imag} */,
  {32'h459bd260, 32'hc46e34e9} /* (12, 27, 31) {real, imag} */,
  {32'hc4d0e6c1, 32'h43093a12} /* (12, 27, 30) {real, imag} */,
  {32'h40c05c70, 32'hc29ec3c2} /* (12, 27, 29) {real, imag} */,
  {32'h425e3e3e, 32'hc38f432e} /* (12, 27, 28) {real, imag} */,
  {32'hc304b16c, 32'h42b98940} /* (12, 27, 27) {real, imag} */,
  {32'hc12303e4, 32'h42b8334e} /* (12, 27, 26) {real, imag} */,
  {32'h418d02ad, 32'hc16de920} /* (12, 27, 25) {real, imag} */,
  {32'hc22239a4, 32'h4330bb64} /* (12, 27, 24) {real, imag} */,
  {32'hc2cd7672, 32'hc25d0d67} /* (12, 27, 23) {real, imag} */,
  {32'h41c774a8, 32'h42a7f2cd} /* (12, 27, 22) {real, imag} */,
  {32'hc19da452, 32'hc03f5640} /* (12, 27, 21) {real, imag} */,
  {32'h430a649e, 32'h42c18f96} /* (12, 27, 20) {real, imag} */,
  {32'hc13c966a, 32'h42e09433} /* (12, 27, 19) {real, imag} */,
  {32'hc1a238c9, 32'hc0911f24} /* (12, 27, 18) {real, imag} */,
  {32'h426d5bd2, 32'h41602e90} /* (12, 27, 17) {real, imag} */,
  {32'h40af9bb4, 32'h00000000} /* (12, 27, 16) {real, imag} */,
  {32'h426d5bd2, 32'hc1602e90} /* (12, 27, 15) {real, imag} */,
  {32'hc1a238c9, 32'h40911f24} /* (12, 27, 14) {real, imag} */,
  {32'hc13c966a, 32'hc2e09433} /* (12, 27, 13) {real, imag} */,
  {32'h430a649e, 32'hc2c18f96} /* (12, 27, 12) {real, imag} */,
  {32'hc19da452, 32'h403f5640} /* (12, 27, 11) {real, imag} */,
  {32'h41c774a8, 32'hc2a7f2cd} /* (12, 27, 10) {real, imag} */,
  {32'hc2cd7672, 32'h425d0d67} /* (12, 27, 9) {real, imag} */,
  {32'hc22239a4, 32'hc330bb64} /* (12, 27, 8) {real, imag} */,
  {32'h418d02ad, 32'h416de920} /* (12, 27, 7) {real, imag} */,
  {32'hc12303e4, 32'hc2b8334e} /* (12, 27, 6) {real, imag} */,
  {32'hc304b16c, 32'hc2b98940} /* (12, 27, 5) {real, imag} */,
  {32'h425e3e3e, 32'h438f432e} /* (12, 27, 4) {real, imag} */,
  {32'h40c05c70, 32'h429ec3c2} /* (12, 27, 3) {real, imag} */,
  {32'hc4d0e6c1, 32'hc3093a12} /* (12, 27, 2) {real, imag} */,
  {32'h459bd260, 32'h446e34e9} /* (12, 27, 1) {real, imag} */,
  {32'h459702f1, 32'h00000000} /* (12, 27, 0) {real, imag} */,
  {32'h4593491a, 32'hc453bc34} /* (12, 26, 31) {real, imag} */,
  {32'hc4da71ea, 32'h4332b962} /* (12, 26, 30) {real, imag} */,
  {32'h4289c3d1, 32'hc2ad5688} /* (12, 26, 29) {real, imag} */,
  {32'h4343d45a, 32'hc200e8e6} /* (12, 26, 28) {real, imag} */,
  {32'hc30dac78, 32'h4319b875} /* (12, 26, 27) {real, imag} */,
  {32'hc2cc7d90, 32'h406ec970} /* (12, 26, 26) {real, imag} */,
  {32'h41aea0ec, 32'hc30dac98} /* (12, 26, 25) {real, imag} */,
  {32'h40ce6e9c, 32'h4324cf60} /* (12, 26, 24) {real, imag} */,
  {32'hc1bbac51, 32'h421ea458} /* (12, 26, 23) {real, imag} */,
  {32'h41ebeb2b, 32'hc2793b0a} /* (12, 26, 22) {real, imag} */,
  {32'h417c2118, 32'h42267fe0} /* (12, 26, 21) {real, imag} */,
  {32'hc2139dd1, 32'h429db610} /* (12, 26, 20) {real, imag} */,
  {32'h421b080c, 32'h427ff571} /* (12, 26, 19) {real, imag} */,
  {32'hc1d63aa4, 32'hc1d968a4} /* (12, 26, 18) {real, imag} */,
  {32'hc1b74629, 32'hc1fba346} /* (12, 26, 17) {real, imag} */,
  {32'hc1bf309b, 32'h00000000} /* (12, 26, 16) {real, imag} */,
  {32'hc1b74629, 32'h41fba346} /* (12, 26, 15) {real, imag} */,
  {32'hc1d63aa4, 32'h41d968a4} /* (12, 26, 14) {real, imag} */,
  {32'h421b080c, 32'hc27ff571} /* (12, 26, 13) {real, imag} */,
  {32'hc2139dd1, 32'hc29db610} /* (12, 26, 12) {real, imag} */,
  {32'h417c2118, 32'hc2267fe0} /* (12, 26, 11) {real, imag} */,
  {32'h41ebeb2b, 32'h42793b0a} /* (12, 26, 10) {real, imag} */,
  {32'hc1bbac51, 32'hc21ea458} /* (12, 26, 9) {real, imag} */,
  {32'h40ce6e9c, 32'hc324cf60} /* (12, 26, 8) {real, imag} */,
  {32'h41aea0ec, 32'h430dac98} /* (12, 26, 7) {real, imag} */,
  {32'hc2cc7d90, 32'hc06ec970} /* (12, 26, 6) {real, imag} */,
  {32'hc30dac78, 32'hc319b875} /* (12, 26, 5) {real, imag} */,
  {32'h4343d45a, 32'h4200e8e6} /* (12, 26, 4) {real, imag} */,
  {32'h4289c3d1, 32'h42ad5688} /* (12, 26, 3) {real, imag} */,
  {32'hc4da71ea, 32'hc332b962} /* (12, 26, 2) {real, imag} */,
  {32'h4593491a, 32'h4453bc34} /* (12, 26, 1) {real, imag} */,
  {32'h458f1f7e, 32'h00000000} /* (12, 26, 0) {real, imag} */,
  {32'h458bb832, 32'hc4336552} /* (12, 25, 31) {real, imag} */,
  {32'hc4d37076, 32'h430ebfca} /* (12, 25, 30) {real, imag} */,
  {32'h41d2d36c, 32'h4215a9f6} /* (12, 25, 29) {real, imag} */,
  {32'h4339a86e, 32'hc28bd2a6} /* (12, 25, 28) {real, imag} */,
  {32'hc2dcfdaa, 32'h4363277d} /* (12, 25, 27) {real, imag} */,
  {32'hc33ebff5, 32'hc2920086} /* (12, 25, 26) {real, imag} */,
  {32'h4252147c, 32'h41fcc7c8} /* (12, 25, 25) {real, imag} */,
  {32'hc2b06a92, 32'h42f03f4d} /* (12, 25, 24) {real, imag} */,
  {32'h427200d2, 32'h3f770700} /* (12, 25, 23) {real, imag} */,
  {32'hc2c8a890, 32'hc3184f53} /* (12, 25, 22) {real, imag} */,
  {32'hc2ac7276, 32'h4234e23a} /* (12, 25, 21) {real, imag} */,
  {32'hc1efe602, 32'h42d40928} /* (12, 25, 20) {real, imag} */,
  {32'h41a31c12, 32'hc229d1e2} /* (12, 25, 19) {real, imag} */,
  {32'h409d0944, 32'h41ad2ea3} /* (12, 25, 18) {real, imag} */,
  {32'h42172d0d, 32'hc29f4a68} /* (12, 25, 17) {real, imag} */,
  {32'h42877a74, 32'h00000000} /* (12, 25, 16) {real, imag} */,
  {32'h42172d0d, 32'h429f4a68} /* (12, 25, 15) {real, imag} */,
  {32'h409d0944, 32'hc1ad2ea3} /* (12, 25, 14) {real, imag} */,
  {32'h41a31c12, 32'h4229d1e2} /* (12, 25, 13) {real, imag} */,
  {32'hc1efe602, 32'hc2d40928} /* (12, 25, 12) {real, imag} */,
  {32'hc2ac7276, 32'hc234e23a} /* (12, 25, 11) {real, imag} */,
  {32'hc2c8a890, 32'h43184f53} /* (12, 25, 10) {real, imag} */,
  {32'h427200d2, 32'hbf770700} /* (12, 25, 9) {real, imag} */,
  {32'hc2b06a92, 32'hc2f03f4d} /* (12, 25, 8) {real, imag} */,
  {32'h4252147c, 32'hc1fcc7c8} /* (12, 25, 7) {real, imag} */,
  {32'hc33ebff5, 32'h42920086} /* (12, 25, 6) {real, imag} */,
  {32'hc2dcfdaa, 32'hc363277d} /* (12, 25, 5) {real, imag} */,
  {32'h4339a86e, 32'h428bd2a6} /* (12, 25, 4) {real, imag} */,
  {32'h41d2d36c, 32'hc215a9f6} /* (12, 25, 3) {real, imag} */,
  {32'hc4d37076, 32'hc30ebfca} /* (12, 25, 2) {real, imag} */,
  {32'h458bb832, 32'h44336552} /* (12, 25, 1) {real, imag} */,
  {32'h457f8be7, 32'h00000000} /* (12, 25, 0) {real, imag} */,
  {32'h457ae782, 32'hc409ac1e} /* (12, 24, 31) {real, imag} */,
  {32'hc4c1f575, 32'h43422592} /* (12, 24, 30) {real, imag} */,
  {32'hc2c71e04, 32'hc230e1b9} /* (12, 24, 29) {real, imag} */,
  {32'h435b5ce8, 32'hc28ca465} /* (12, 24, 28) {real, imag} */,
  {32'hc2a79677, 32'h43489e52} /* (12, 24, 27) {real, imag} */,
  {32'hc3179ed8, 32'hc27423a0} /* (12, 24, 26) {real, imag} */,
  {32'h42b7459c, 32'hc1f71943} /* (12, 24, 25) {real, imag} */,
  {32'hc2939b62, 32'h434679e2} /* (12, 24, 24) {real, imag} */,
  {32'h42b55f1a, 32'h426973be} /* (12, 24, 23) {real, imag} */,
  {32'h41b78d62, 32'hc31e7976} /* (12, 24, 22) {real, imag} */,
  {32'hc215b72b, 32'h42ab42c7} /* (12, 24, 21) {real, imag} */,
  {32'h417cfa28, 32'hc1f297b4} /* (12, 24, 20) {real, imag} */,
  {32'hc0c7a8a0, 32'hc2abc475} /* (12, 24, 19) {real, imag} */,
  {32'h41d0f8c3, 32'hc19b271e} /* (12, 24, 18) {real, imag} */,
  {32'h40bab9e4, 32'h422bf532} /* (12, 24, 17) {real, imag} */,
  {32'h3ff5ba20, 32'h00000000} /* (12, 24, 16) {real, imag} */,
  {32'h40bab9e4, 32'hc22bf532} /* (12, 24, 15) {real, imag} */,
  {32'h41d0f8c3, 32'h419b271e} /* (12, 24, 14) {real, imag} */,
  {32'hc0c7a8a0, 32'h42abc475} /* (12, 24, 13) {real, imag} */,
  {32'h417cfa28, 32'h41f297b4} /* (12, 24, 12) {real, imag} */,
  {32'hc215b72b, 32'hc2ab42c7} /* (12, 24, 11) {real, imag} */,
  {32'h41b78d62, 32'h431e7976} /* (12, 24, 10) {real, imag} */,
  {32'h42b55f1a, 32'hc26973be} /* (12, 24, 9) {real, imag} */,
  {32'hc2939b62, 32'hc34679e2} /* (12, 24, 8) {real, imag} */,
  {32'h42b7459c, 32'h41f71943} /* (12, 24, 7) {real, imag} */,
  {32'hc3179ed8, 32'h427423a0} /* (12, 24, 6) {real, imag} */,
  {32'hc2a79677, 32'hc3489e52} /* (12, 24, 5) {real, imag} */,
  {32'h435b5ce8, 32'h428ca465} /* (12, 24, 4) {real, imag} */,
  {32'hc2c71e04, 32'h4230e1b9} /* (12, 24, 3) {real, imag} */,
  {32'hc4c1f575, 32'hc3422592} /* (12, 24, 2) {real, imag} */,
  {32'h457ae782, 32'h4409ac1e} /* (12, 24, 1) {real, imag} */,
  {32'h45588330, 32'h00000000} /* (12, 24, 0) {real, imag} */,
  {32'h454cdd4d, 32'hc3ff7483} /* (12, 23, 31) {real, imag} */,
  {32'hc4973298, 32'h432cbfa7} /* (12, 23, 30) {real, imag} */,
  {32'hc2f17597, 32'hc2062a82} /* (12, 23, 29) {real, imag} */,
  {32'h4325dbd5, 32'hc333a8cf} /* (12, 23, 28) {real, imag} */,
  {32'hc3681963, 32'h42877658} /* (12, 23, 27) {real, imag} */,
  {32'hc24aa5cb, 32'h418644a1} /* (12, 23, 26) {real, imag} */,
  {32'hc0d84ca4, 32'hc1e49194} /* (12, 23, 25) {real, imag} */,
  {32'hc102901e, 32'h426b23fe} /* (12, 23, 24) {real, imag} */,
  {32'hc29ea9d4, 32'h428acc25} /* (12, 23, 23) {real, imag} */,
  {32'h420f9cdf, 32'h42932a49} /* (12, 23, 22) {real, imag} */,
  {32'h4277d3e5, 32'h4262c04a} /* (12, 23, 21) {real, imag} */,
  {32'hc262c994, 32'h42098d84} /* (12, 23, 20) {real, imag} */,
  {32'h4252d5ba, 32'h40ee4440} /* (12, 23, 19) {real, imag} */,
  {32'hc093d6a0, 32'hc07b7bb0} /* (12, 23, 18) {real, imag} */,
  {32'h416980f2, 32'hc284cd3e} /* (12, 23, 17) {real, imag} */,
  {32'hc21c6080, 32'h00000000} /* (12, 23, 16) {real, imag} */,
  {32'h416980f2, 32'h4284cd3e} /* (12, 23, 15) {real, imag} */,
  {32'hc093d6a0, 32'h407b7bb0} /* (12, 23, 14) {real, imag} */,
  {32'h4252d5ba, 32'hc0ee4440} /* (12, 23, 13) {real, imag} */,
  {32'hc262c994, 32'hc2098d84} /* (12, 23, 12) {real, imag} */,
  {32'h4277d3e5, 32'hc262c04a} /* (12, 23, 11) {real, imag} */,
  {32'h420f9cdf, 32'hc2932a49} /* (12, 23, 10) {real, imag} */,
  {32'hc29ea9d4, 32'hc28acc25} /* (12, 23, 9) {real, imag} */,
  {32'hc102901e, 32'hc26b23fe} /* (12, 23, 8) {real, imag} */,
  {32'hc0d84ca4, 32'h41e49194} /* (12, 23, 7) {real, imag} */,
  {32'hc24aa5cb, 32'hc18644a1} /* (12, 23, 6) {real, imag} */,
  {32'hc3681963, 32'hc2877658} /* (12, 23, 5) {real, imag} */,
  {32'h4325dbd5, 32'h4333a8cf} /* (12, 23, 4) {real, imag} */,
  {32'hc2f17597, 32'h42062a82} /* (12, 23, 3) {real, imag} */,
  {32'hc4973298, 32'hc32cbfa7} /* (12, 23, 2) {real, imag} */,
  {32'h454cdd4d, 32'h43ff7483} /* (12, 23, 1) {real, imag} */,
  {32'h45284369, 32'h00000000} /* (12, 23, 0) {real, imag} */,
  {32'h4515661e, 32'hc39c888f} /* (12, 22, 31) {real, imag} */,
  {32'hc44fcd15, 32'h4354b89e} /* (12, 22, 30) {real, imag} */,
  {32'hc257e2c2, 32'hc1bebde2} /* (12, 22, 29) {real, imag} */,
  {32'h43ac0825, 32'hc33c6a4e} /* (12, 22, 28) {real, imag} */,
  {32'hc38e7d5a, 32'h4368e7a8} /* (12, 22, 27) {real, imag} */,
  {32'hc320d61c, 32'hc2736e6d} /* (12, 22, 26) {real, imag} */,
  {32'h430e42ea, 32'h40ea7be8} /* (12, 22, 25) {real, imag} */,
  {32'hc30e6251, 32'hc119bc2c} /* (12, 22, 24) {real, imag} */,
  {32'hc2c93aaa, 32'h42c9fedf} /* (12, 22, 23) {real, imag} */,
  {32'h42b3f2d9, 32'h41ab91e9} /* (12, 22, 22) {real, imag} */,
  {32'hc2a3ec6a, 32'h41bd98b4} /* (12, 22, 21) {real, imag} */,
  {32'hc23dccf2, 32'h421c17f5} /* (12, 22, 20) {real, imag} */,
  {32'h40146460, 32'h418d6ebf} /* (12, 22, 19) {real, imag} */,
  {32'h420bde1c, 32'hc128b978} /* (12, 22, 18) {real, imag} */,
  {32'h42b92176, 32'h42191198} /* (12, 22, 17) {real, imag} */,
  {32'hc2fd70d2, 32'h00000000} /* (12, 22, 16) {real, imag} */,
  {32'h42b92176, 32'hc2191198} /* (12, 22, 15) {real, imag} */,
  {32'h420bde1c, 32'h4128b978} /* (12, 22, 14) {real, imag} */,
  {32'h40146460, 32'hc18d6ebf} /* (12, 22, 13) {real, imag} */,
  {32'hc23dccf2, 32'hc21c17f5} /* (12, 22, 12) {real, imag} */,
  {32'hc2a3ec6a, 32'hc1bd98b4} /* (12, 22, 11) {real, imag} */,
  {32'h42b3f2d9, 32'hc1ab91e9} /* (12, 22, 10) {real, imag} */,
  {32'hc2c93aaa, 32'hc2c9fedf} /* (12, 22, 9) {real, imag} */,
  {32'hc30e6251, 32'h4119bc2c} /* (12, 22, 8) {real, imag} */,
  {32'h430e42ea, 32'hc0ea7be8} /* (12, 22, 7) {real, imag} */,
  {32'hc320d61c, 32'h42736e6d} /* (12, 22, 6) {real, imag} */,
  {32'hc38e7d5a, 32'hc368e7a8} /* (12, 22, 5) {real, imag} */,
  {32'h43ac0825, 32'h433c6a4e} /* (12, 22, 4) {real, imag} */,
  {32'hc257e2c2, 32'h41bebde2} /* (12, 22, 3) {real, imag} */,
  {32'hc44fcd15, 32'hc354b89e} /* (12, 22, 2) {real, imag} */,
  {32'h4515661e, 32'h439c888f} /* (12, 22, 1) {real, imag} */,
  {32'h44e815af, 32'h00000000} /* (12, 22, 0) {real, imag} */,
  {32'h443c8e7c, 32'h40bee100} /* (12, 21, 31) {real, imag} */,
  {32'hc378b440, 32'h414d0a60} /* (12, 21, 30) {real, imag} */,
  {32'hc23b3ecf, 32'hc13efeae} /* (12, 21, 29) {real, imag} */,
  {32'h433f8de4, 32'hc17ec510} /* (12, 21, 28) {real, imag} */,
  {32'hc3260b0a, 32'h42e31250} /* (12, 21, 27) {real, imag} */,
  {32'hc2ab5b1e, 32'h4141025e} /* (12, 21, 26) {real, imag} */,
  {32'h42135774, 32'hc1941bd4} /* (12, 21, 25) {real, imag} */,
  {32'hc2cbf3a8, 32'h404ec0bc} /* (12, 21, 24) {real, imag} */,
  {32'h4272d1a5, 32'h40c846fa} /* (12, 21, 23) {real, imag} */,
  {32'hc1cbfd5a, 32'hc2c2c8df} /* (12, 21, 22) {real, imag} */,
  {32'hc2c699ea, 32'h41aa8fe2} /* (12, 21, 21) {real, imag} */,
  {32'hc2347020, 32'hc2774280} /* (12, 21, 20) {real, imag} */,
  {32'hc1b29244, 32'h4198b10b} /* (12, 21, 19) {real, imag} */,
  {32'hc0b47ae4, 32'h41c30518} /* (12, 21, 18) {real, imag} */,
  {32'hc1ff46e4, 32'h4194ad3a} /* (12, 21, 17) {real, imag} */,
  {32'h4302e420, 32'h00000000} /* (12, 21, 16) {real, imag} */,
  {32'hc1ff46e4, 32'hc194ad3a} /* (12, 21, 15) {real, imag} */,
  {32'hc0b47ae4, 32'hc1c30518} /* (12, 21, 14) {real, imag} */,
  {32'hc1b29244, 32'hc198b10b} /* (12, 21, 13) {real, imag} */,
  {32'hc2347020, 32'h42774280} /* (12, 21, 12) {real, imag} */,
  {32'hc2c699ea, 32'hc1aa8fe2} /* (12, 21, 11) {real, imag} */,
  {32'hc1cbfd5a, 32'h42c2c8df} /* (12, 21, 10) {real, imag} */,
  {32'h4272d1a5, 32'hc0c846fa} /* (12, 21, 9) {real, imag} */,
  {32'hc2cbf3a8, 32'hc04ec0bc} /* (12, 21, 8) {real, imag} */,
  {32'h42135774, 32'h41941bd4} /* (12, 21, 7) {real, imag} */,
  {32'hc2ab5b1e, 32'hc141025e} /* (12, 21, 6) {real, imag} */,
  {32'hc3260b0a, 32'hc2e31250} /* (12, 21, 5) {real, imag} */,
  {32'h433f8de4, 32'h417ec510} /* (12, 21, 4) {real, imag} */,
  {32'hc23b3ecf, 32'h413efeae} /* (12, 21, 3) {real, imag} */,
  {32'hc378b440, 32'hc14d0a60} /* (12, 21, 2) {real, imag} */,
  {32'h443c8e7c, 32'hc0bee100} /* (12, 21, 1) {real, imag} */,
  {32'h442db1ad, 32'h00000000} /* (12, 21, 0) {real, imag} */,
  {32'hc49515b8, 32'h435316a4} /* (12, 20, 31) {real, imag} */,
  {32'h441ac181, 32'hc313305f} /* (12, 20, 30) {real, imag} */,
  {32'hc300b7b5, 32'h4191908a} /* (12, 20, 29) {real, imag} */,
  {32'hc253da1a, 32'h433ca5da} /* (12, 20, 28) {real, imag} */,
  {32'h4353ddca, 32'hc2208e58} /* (12, 20, 27) {real, imag} */,
  {32'h41fcd5d8, 32'h4197b207} /* (12, 20, 26) {real, imag} */,
  {32'hc28ad458, 32'hc1052148} /* (12, 20, 25) {real, imag} */,
  {32'h42c2d10c, 32'hc1d85544} /* (12, 20, 24) {real, imag} */,
  {32'h42725482, 32'hc20b3e0e} /* (12, 20, 23) {real, imag} */,
  {32'hc2cd1afc, 32'h4273d632} /* (12, 20, 22) {real, imag} */,
  {32'h42c0dba5, 32'hc1761f44} /* (12, 20, 21) {real, imag} */,
  {32'hc142fd6c, 32'hc2a4b0c2} /* (12, 20, 20) {real, imag} */,
  {32'h41ca90ad, 32'hc268e476} /* (12, 20, 19) {real, imag} */,
  {32'hc2ae779d, 32'h41a2333a} /* (12, 20, 18) {real, imag} */,
  {32'h4234cda2, 32'hc2d85af7} /* (12, 20, 17) {real, imag} */,
  {32'hc1980dc2, 32'h00000000} /* (12, 20, 16) {real, imag} */,
  {32'h4234cda2, 32'h42d85af7} /* (12, 20, 15) {real, imag} */,
  {32'hc2ae779d, 32'hc1a2333a} /* (12, 20, 14) {real, imag} */,
  {32'h41ca90ad, 32'h4268e476} /* (12, 20, 13) {real, imag} */,
  {32'hc142fd6c, 32'h42a4b0c2} /* (12, 20, 12) {real, imag} */,
  {32'h42c0dba5, 32'h41761f44} /* (12, 20, 11) {real, imag} */,
  {32'hc2cd1afc, 32'hc273d632} /* (12, 20, 10) {real, imag} */,
  {32'h42725482, 32'h420b3e0e} /* (12, 20, 9) {real, imag} */,
  {32'h42c2d10c, 32'h41d85544} /* (12, 20, 8) {real, imag} */,
  {32'hc28ad458, 32'h41052148} /* (12, 20, 7) {real, imag} */,
  {32'h41fcd5d8, 32'hc197b207} /* (12, 20, 6) {real, imag} */,
  {32'h4353ddca, 32'h42208e58} /* (12, 20, 5) {real, imag} */,
  {32'hc253da1a, 32'hc33ca5da} /* (12, 20, 4) {real, imag} */,
  {32'hc300b7b5, 32'hc191908a} /* (12, 20, 3) {real, imag} */,
  {32'h441ac181, 32'h4313305f} /* (12, 20, 2) {real, imag} */,
  {32'hc49515b8, 32'hc35316a4} /* (12, 20, 1) {real, imag} */,
  {32'hc45728fe, 32'h00000000} /* (12, 20, 0) {real, imag} */,
  {32'hc514c6b1, 32'h43847d78} /* (12, 19, 31) {real, imag} */,
  {32'h4485a3ec, 32'hc36a2a15} /* (12, 19, 30) {real, imag} */,
  {32'hc2d16014, 32'h41340602} /* (12, 19, 29) {real, imag} */,
  {32'hc2cac844, 32'h426ade06} /* (12, 19, 28) {real, imag} */,
  {32'h4333ff7b, 32'h41c0d4ae} /* (12, 19, 27) {real, imag} */,
  {32'hc28cda5c, 32'hc200ce83} /* (12, 19, 26) {real, imag} */,
  {32'hc2bca94e, 32'h428424b2} /* (12, 19, 25) {real, imag} */,
  {32'h42defd2b, 32'hc33dc0e7} /* (12, 19, 24) {real, imag} */,
  {32'h41c70835, 32'hc21ea360} /* (12, 19, 23) {real, imag} */,
  {32'hc17d7fd8, 32'hc2e02748} /* (12, 19, 22) {real, imag} */,
  {32'h42a67cf8, 32'hc299350d} /* (12, 19, 21) {real, imag} */,
  {32'h428180c0, 32'h41915414} /* (12, 19, 20) {real, imag} */,
  {32'hc1536a84, 32'h420fc56a} /* (12, 19, 19) {real, imag} */,
  {32'hc2e3cdeb, 32'hc2d4a0e6} /* (12, 19, 18) {real, imag} */,
  {32'hc27b285f, 32'hc149c9c8} /* (12, 19, 17) {real, imag} */,
  {32'hc0e76e0c, 32'h00000000} /* (12, 19, 16) {real, imag} */,
  {32'hc27b285f, 32'h4149c9c8} /* (12, 19, 15) {real, imag} */,
  {32'hc2e3cdeb, 32'h42d4a0e6} /* (12, 19, 14) {real, imag} */,
  {32'hc1536a84, 32'hc20fc56a} /* (12, 19, 13) {real, imag} */,
  {32'h428180c0, 32'hc1915414} /* (12, 19, 12) {real, imag} */,
  {32'h42a67cf8, 32'h4299350d} /* (12, 19, 11) {real, imag} */,
  {32'hc17d7fd8, 32'h42e02748} /* (12, 19, 10) {real, imag} */,
  {32'h41c70835, 32'h421ea360} /* (12, 19, 9) {real, imag} */,
  {32'h42defd2b, 32'h433dc0e7} /* (12, 19, 8) {real, imag} */,
  {32'hc2bca94e, 32'hc28424b2} /* (12, 19, 7) {real, imag} */,
  {32'hc28cda5c, 32'h4200ce83} /* (12, 19, 6) {real, imag} */,
  {32'h4333ff7b, 32'hc1c0d4ae} /* (12, 19, 5) {real, imag} */,
  {32'hc2cac844, 32'hc26ade06} /* (12, 19, 4) {real, imag} */,
  {32'hc2d16014, 32'hc1340602} /* (12, 19, 3) {real, imag} */,
  {32'h4485a3ec, 32'h436a2a15} /* (12, 19, 2) {real, imag} */,
  {32'hc514c6b1, 32'hc3847d78} /* (12, 19, 1) {real, imag} */,
  {32'hc4def6e4, 32'h00000000} /* (12, 19, 0) {real, imag} */,
  {32'hc5490edd, 32'h43e8c616} /* (12, 18, 31) {real, imag} */,
  {32'h44a4e7e4, 32'hc38328b1} /* (12, 18, 30) {real, imag} */,
  {32'hc1980178, 32'h4161b008} /* (12, 18, 29) {real, imag} */,
  {32'hc293b25c, 32'h4309b374} /* (12, 18, 28) {real, imag} */,
  {32'h43a9d41c, 32'hc3197dfc} /* (12, 18, 27) {real, imag} */,
  {32'hc275d68c, 32'h41b87a34} /* (12, 18, 26) {real, imag} */,
  {32'h418bbbf6, 32'hc1eacdc6} /* (12, 18, 25) {real, imag} */,
  {32'h41d70136, 32'hc2cb5eaa} /* (12, 18, 24) {real, imag} */,
  {32'h42e6aa66, 32'h42363788} /* (12, 18, 23) {real, imag} */,
  {32'hc2a42020, 32'h428d8a4d} /* (12, 18, 22) {real, imag} */,
  {32'hc20fdf4f, 32'hc29e487e} /* (12, 18, 21) {real, imag} */,
  {32'hc218580a, 32'h42855ced} /* (12, 18, 20) {real, imag} */,
  {32'h41945cee, 32'h430a6f55} /* (12, 18, 19) {real, imag} */,
  {32'h419e6448, 32'hc2c93f72} /* (12, 18, 18) {real, imag} */,
  {32'hc22a10cc, 32'h42507e48} /* (12, 18, 17) {real, imag} */,
  {32'h42926c80, 32'h00000000} /* (12, 18, 16) {real, imag} */,
  {32'hc22a10cc, 32'hc2507e48} /* (12, 18, 15) {real, imag} */,
  {32'h419e6448, 32'h42c93f72} /* (12, 18, 14) {real, imag} */,
  {32'h41945cee, 32'hc30a6f55} /* (12, 18, 13) {real, imag} */,
  {32'hc218580a, 32'hc2855ced} /* (12, 18, 12) {real, imag} */,
  {32'hc20fdf4f, 32'h429e487e} /* (12, 18, 11) {real, imag} */,
  {32'hc2a42020, 32'hc28d8a4d} /* (12, 18, 10) {real, imag} */,
  {32'h42e6aa66, 32'hc2363788} /* (12, 18, 9) {real, imag} */,
  {32'h41d70136, 32'h42cb5eaa} /* (12, 18, 8) {real, imag} */,
  {32'h418bbbf6, 32'h41eacdc6} /* (12, 18, 7) {real, imag} */,
  {32'hc275d68c, 32'hc1b87a34} /* (12, 18, 6) {real, imag} */,
  {32'h43a9d41c, 32'h43197dfc} /* (12, 18, 5) {real, imag} */,
  {32'hc293b25c, 32'hc309b374} /* (12, 18, 4) {real, imag} */,
  {32'hc1980178, 32'hc161b008} /* (12, 18, 3) {real, imag} */,
  {32'h44a4e7e4, 32'h438328b1} /* (12, 18, 2) {real, imag} */,
  {32'hc5490edd, 32'hc3e8c616} /* (12, 18, 1) {real, imag} */,
  {32'hc51fd213, 32'h00000000} /* (12, 18, 0) {real, imag} */,
  {32'hc56c6054, 32'h43fe8a6d} /* (12, 17, 31) {real, imag} */,
  {32'h44bbf0e9, 32'hc36fd60a} /* (12, 17, 30) {real, imag} */,
  {32'h42e237ab, 32'h413c84c2} /* (12, 17, 29) {real, imag} */,
  {32'h421f3cfc, 32'h42a1cdb6} /* (12, 17, 28) {real, imag} */,
  {32'h43ac8af7, 32'hc2cc8709} /* (12, 17, 27) {real, imag} */,
  {32'h41d007e4, 32'hc2ac40b0} /* (12, 17, 26) {real, imag} */,
  {32'hc2e7a44d, 32'h40cf8860} /* (12, 17, 25) {real, imag} */,
  {32'hbfc53a00, 32'h419feaae} /* (12, 17, 24) {real, imag} */,
  {32'hc2b47806, 32'h42d75d19} /* (12, 17, 23) {real, imag} */,
  {32'hc22cc61e, 32'hc1b17276} /* (12, 17, 22) {real, imag} */,
  {32'h428a28ce, 32'h4165559a} /* (12, 17, 21) {real, imag} */,
  {32'hc24ee68b, 32'hc15b3ed6} /* (12, 17, 20) {real, imag} */,
  {32'h4211c668, 32'hc26d9096} /* (12, 17, 19) {real, imag} */,
  {32'hc23e7b43, 32'hc2a870c7} /* (12, 17, 18) {real, imag} */,
  {32'hc23656be, 32'h41e4b494} /* (12, 17, 17) {real, imag} */,
  {32'hc2307148, 32'h00000000} /* (12, 17, 16) {real, imag} */,
  {32'hc23656be, 32'hc1e4b494} /* (12, 17, 15) {real, imag} */,
  {32'hc23e7b43, 32'h42a870c7} /* (12, 17, 14) {real, imag} */,
  {32'h4211c668, 32'h426d9096} /* (12, 17, 13) {real, imag} */,
  {32'hc24ee68b, 32'h415b3ed6} /* (12, 17, 12) {real, imag} */,
  {32'h428a28ce, 32'hc165559a} /* (12, 17, 11) {real, imag} */,
  {32'hc22cc61e, 32'h41b17276} /* (12, 17, 10) {real, imag} */,
  {32'hc2b47806, 32'hc2d75d19} /* (12, 17, 9) {real, imag} */,
  {32'hbfc53a00, 32'hc19feaae} /* (12, 17, 8) {real, imag} */,
  {32'hc2e7a44d, 32'hc0cf8860} /* (12, 17, 7) {real, imag} */,
  {32'h41d007e4, 32'h42ac40b0} /* (12, 17, 6) {real, imag} */,
  {32'h43ac8af7, 32'h42cc8709} /* (12, 17, 5) {real, imag} */,
  {32'h421f3cfc, 32'hc2a1cdb6} /* (12, 17, 4) {real, imag} */,
  {32'h42e237ab, 32'hc13c84c2} /* (12, 17, 3) {real, imag} */,
  {32'h44bbf0e9, 32'h436fd60a} /* (12, 17, 2) {real, imag} */,
  {32'hc56c6054, 32'hc3fe8a6d} /* (12, 17, 1) {real, imag} */,
  {32'hc536137e, 32'h00000000} /* (12, 17, 0) {real, imag} */,
  {32'hc57fd375, 32'h4404760e} /* (12, 16, 31) {real, imag} */,
  {32'h44c2a904, 32'hc35c3a96} /* (12, 16, 30) {real, imag} */,
  {32'h42573853, 32'hc2c91d08} /* (12, 16, 29) {real, imag} */,
  {32'hc36569f0, 32'h42cb0b0a} /* (12, 16, 28) {real, imag} */,
  {32'h43817905, 32'h425700b0} /* (12, 16, 27) {real, imag} */,
  {32'hc290e458, 32'hc19a5346} /* (12, 16, 26) {real, imag} */,
  {32'hc2857760, 32'hc15a2ecc} /* (12, 16, 25) {real, imag} */,
  {32'h42bfb4e1, 32'h4218e2fc} /* (12, 16, 24) {real, imag} */,
  {32'hc2b810b0, 32'hc2766848} /* (12, 16, 23) {real, imag} */,
  {32'hc29b5d4c, 32'hc24db47b} /* (12, 16, 22) {real, imag} */,
  {32'hc23713b4, 32'hc2c1a592} /* (12, 16, 21) {real, imag} */,
  {32'h421a701d, 32'hc2905dbb} /* (12, 16, 20) {real, imag} */,
  {32'hc1f75645, 32'h404c8330} /* (12, 16, 19) {real, imag} */,
  {32'h426fee55, 32'hc1f96acc} /* (12, 16, 18) {real, imag} */,
  {32'hc1c1a800, 32'hc25aaa66} /* (12, 16, 17) {real, imag} */,
  {32'h4290c604, 32'h00000000} /* (12, 16, 16) {real, imag} */,
  {32'hc1c1a800, 32'h425aaa66} /* (12, 16, 15) {real, imag} */,
  {32'h426fee55, 32'h41f96acc} /* (12, 16, 14) {real, imag} */,
  {32'hc1f75645, 32'hc04c8330} /* (12, 16, 13) {real, imag} */,
  {32'h421a701d, 32'h42905dbb} /* (12, 16, 12) {real, imag} */,
  {32'hc23713b4, 32'h42c1a592} /* (12, 16, 11) {real, imag} */,
  {32'hc29b5d4c, 32'h424db47b} /* (12, 16, 10) {real, imag} */,
  {32'hc2b810b0, 32'h42766848} /* (12, 16, 9) {real, imag} */,
  {32'h42bfb4e1, 32'hc218e2fc} /* (12, 16, 8) {real, imag} */,
  {32'hc2857760, 32'h415a2ecc} /* (12, 16, 7) {real, imag} */,
  {32'hc290e458, 32'h419a5346} /* (12, 16, 6) {real, imag} */,
  {32'h43817905, 32'hc25700b0} /* (12, 16, 5) {real, imag} */,
  {32'hc36569f0, 32'hc2cb0b0a} /* (12, 16, 4) {real, imag} */,
  {32'h42573853, 32'h42c91d08} /* (12, 16, 3) {real, imag} */,
  {32'h44c2a904, 32'h435c3a96} /* (12, 16, 2) {real, imag} */,
  {32'hc57fd375, 32'hc404760e} /* (12, 16, 1) {real, imag} */,
  {32'hc53d5b76, 32'h00000000} /* (12, 16, 0) {real, imag} */,
  {32'hc58030aa, 32'h43e639d3} /* (12, 15, 31) {real, imag} */,
  {32'h44b6392b, 32'hc335350a} /* (12, 15, 30) {real, imag} */,
  {32'h42767e06, 32'hc25fbce4} /* (12, 15, 29) {real, imag} */,
  {32'hc36a1985, 32'h42a2028a} /* (12, 15, 28) {real, imag} */,
  {32'h42be9265, 32'hc2a35a27} /* (12, 15, 27) {real, imag} */,
  {32'hc293c2a6, 32'hc295787a} /* (12, 15, 26) {real, imag} */,
  {32'hc24b2dfe, 32'hc2c0d77c} /* (12, 15, 25) {real, imag} */,
  {32'hc22d1730, 32'h4125f00a} /* (12, 15, 24) {real, imag} */,
  {32'hc2b77566, 32'h423d9286} /* (12, 15, 23) {real, imag} */,
  {32'hc25fe576, 32'h41fc8c62} /* (12, 15, 22) {real, imag} */,
  {32'h41859a1a, 32'hc19f4e99} /* (12, 15, 21) {real, imag} */,
  {32'hc184d00e, 32'hc2829c26} /* (12, 15, 20) {real, imag} */,
  {32'h41313ac0, 32'hc285cb51} /* (12, 15, 19) {real, imag} */,
  {32'h410f8ea0, 32'hc1d1c81d} /* (12, 15, 18) {real, imag} */,
  {32'hc25c7326, 32'hc1234bcf} /* (12, 15, 17) {real, imag} */,
  {32'hc2b7e92a, 32'h00000000} /* (12, 15, 16) {real, imag} */,
  {32'hc25c7326, 32'h41234bcf} /* (12, 15, 15) {real, imag} */,
  {32'h410f8ea0, 32'h41d1c81d} /* (12, 15, 14) {real, imag} */,
  {32'h41313ac0, 32'h4285cb51} /* (12, 15, 13) {real, imag} */,
  {32'hc184d00e, 32'h42829c26} /* (12, 15, 12) {real, imag} */,
  {32'h41859a1a, 32'h419f4e99} /* (12, 15, 11) {real, imag} */,
  {32'hc25fe576, 32'hc1fc8c62} /* (12, 15, 10) {real, imag} */,
  {32'hc2b77566, 32'hc23d9286} /* (12, 15, 9) {real, imag} */,
  {32'hc22d1730, 32'hc125f00a} /* (12, 15, 8) {real, imag} */,
  {32'hc24b2dfe, 32'h42c0d77c} /* (12, 15, 7) {real, imag} */,
  {32'hc293c2a6, 32'h4295787a} /* (12, 15, 6) {real, imag} */,
  {32'h42be9265, 32'h42a35a27} /* (12, 15, 5) {real, imag} */,
  {32'hc36a1985, 32'hc2a2028a} /* (12, 15, 4) {real, imag} */,
  {32'h42767e06, 32'h425fbce4} /* (12, 15, 3) {real, imag} */,
  {32'h44b6392b, 32'h4335350a} /* (12, 15, 2) {real, imag} */,
  {32'hc58030aa, 32'hc3e639d3} /* (12, 15, 1) {real, imag} */,
  {32'hc544275e, 32'h00000000} /* (12, 15, 0) {real, imag} */,
  {32'hc576f82f, 32'h43bf44c2} /* (12, 14, 31) {real, imag} */,
  {32'h44a846ec, 32'hc37a9ce6} /* (12, 14, 30) {real, imag} */,
  {32'h419b9f08, 32'h42ae4e8a} /* (12, 14, 29) {real, imag} */,
  {32'hc3879cbd, 32'h43207894} /* (12, 14, 28) {real, imag} */,
  {32'hc2b37a30, 32'hc333d408} /* (12, 14, 27) {real, imag} */,
  {32'hc27dc5d6, 32'hc346b52c} /* (12, 14, 26) {real, imag} */,
  {32'hc2266de1, 32'h41bc3352} /* (12, 14, 25) {real, imag} */,
  {32'h41ffda32, 32'hc11c4fe4} /* (12, 14, 24) {real, imag} */,
  {32'hc09cbc88, 32'h4107be56} /* (12, 14, 23) {real, imag} */,
  {32'hc2925afc, 32'hc26ff2be} /* (12, 14, 22) {real, imag} */,
  {32'h42531925, 32'hc3102bcf} /* (12, 14, 21) {real, imag} */,
  {32'hc10438be, 32'hc1a1723d} /* (12, 14, 20) {real, imag} */,
  {32'h42826a16, 32'h41d4ef00} /* (12, 14, 19) {real, imag} */,
  {32'hc21eac3e, 32'hc24b4029} /* (12, 14, 18) {real, imag} */,
  {32'hc0014758, 32'h41835d1c} /* (12, 14, 17) {real, imag} */,
  {32'h41b737d6, 32'h00000000} /* (12, 14, 16) {real, imag} */,
  {32'hc0014758, 32'hc1835d1c} /* (12, 14, 15) {real, imag} */,
  {32'hc21eac3e, 32'h424b4029} /* (12, 14, 14) {real, imag} */,
  {32'h42826a16, 32'hc1d4ef00} /* (12, 14, 13) {real, imag} */,
  {32'hc10438be, 32'h41a1723d} /* (12, 14, 12) {real, imag} */,
  {32'h42531925, 32'h43102bcf} /* (12, 14, 11) {real, imag} */,
  {32'hc2925afc, 32'h426ff2be} /* (12, 14, 10) {real, imag} */,
  {32'hc09cbc88, 32'hc107be56} /* (12, 14, 9) {real, imag} */,
  {32'h41ffda32, 32'h411c4fe4} /* (12, 14, 8) {real, imag} */,
  {32'hc2266de1, 32'hc1bc3352} /* (12, 14, 7) {real, imag} */,
  {32'hc27dc5d6, 32'h4346b52c} /* (12, 14, 6) {real, imag} */,
  {32'hc2b37a30, 32'h4333d408} /* (12, 14, 5) {real, imag} */,
  {32'hc3879cbd, 32'hc3207894} /* (12, 14, 4) {real, imag} */,
  {32'h419b9f08, 32'hc2ae4e8a} /* (12, 14, 3) {real, imag} */,
  {32'h44a846ec, 32'h437a9ce6} /* (12, 14, 2) {real, imag} */,
  {32'hc576f82f, 32'hc3bf44c2} /* (12, 14, 1) {real, imag} */,
  {32'hc535be81, 32'h00000000} /* (12, 14, 0) {real, imag} */,
  {32'hc558e24b, 32'h439704c8} /* (12, 13, 31) {real, imag} */,
  {32'h448f9cb0, 32'hc344e0df} /* (12, 13, 30) {real, imag} */,
  {32'hc301c3a6, 32'h41eae699} /* (12, 13, 29) {real, imag} */,
  {32'hc345344a, 32'h4367fa72} /* (12, 13, 28) {real, imag} */,
  {32'h43713c95, 32'hc2e06428} /* (12, 13, 27) {real, imag} */,
  {32'h4239dee5, 32'hc2fc5c32} /* (12, 13, 26) {real, imag} */,
  {32'h41827e4e, 32'hc207396a} /* (12, 13, 25) {real, imag} */,
  {32'hc16adc30, 32'hc25f9244} /* (12, 13, 24) {real, imag} */,
  {32'h42582a54, 32'hc0ecad20} /* (12, 13, 23) {real, imag} */,
  {32'hc200a19a, 32'h3fd62c00} /* (12, 13, 22) {real, imag} */,
  {32'h4337cc58, 32'hc301aa15} /* (12, 13, 21) {real, imag} */,
  {32'h42268746, 32'hc1d42e60} /* (12, 13, 20) {real, imag} */,
  {32'hc2815c3c, 32'h420c3a6a} /* (12, 13, 19) {real, imag} */,
  {32'h4162c268, 32'hc0928f40} /* (12, 13, 18) {real, imag} */,
  {32'hc284a976, 32'hc1c4f144} /* (12, 13, 17) {real, imag} */,
  {32'hc10738fe, 32'h00000000} /* (12, 13, 16) {real, imag} */,
  {32'hc284a976, 32'h41c4f144} /* (12, 13, 15) {real, imag} */,
  {32'h4162c268, 32'h40928f40} /* (12, 13, 14) {real, imag} */,
  {32'hc2815c3c, 32'hc20c3a6a} /* (12, 13, 13) {real, imag} */,
  {32'h42268746, 32'h41d42e60} /* (12, 13, 12) {real, imag} */,
  {32'h4337cc58, 32'h4301aa15} /* (12, 13, 11) {real, imag} */,
  {32'hc200a19a, 32'hbfd62c00} /* (12, 13, 10) {real, imag} */,
  {32'h42582a54, 32'h40ecad20} /* (12, 13, 9) {real, imag} */,
  {32'hc16adc30, 32'h425f9244} /* (12, 13, 8) {real, imag} */,
  {32'h41827e4e, 32'h4207396a} /* (12, 13, 7) {real, imag} */,
  {32'h4239dee5, 32'h42fc5c32} /* (12, 13, 6) {real, imag} */,
  {32'h43713c95, 32'h42e06428} /* (12, 13, 5) {real, imag} */,
  {32'hc345344a, 32'hc367fa72} /* (12, 13, 4) {real, imag} */,
  {32'hc301c3a6, 32'hc1eae699} /* (12, 13, 3) {real, imag} */,
  {32'h448f9cb0, 32'h4344e0df} /* (12, 13, 2) {real, imag} */,
  {32'hc558e24b, 32'hc39704c8} /* (12, 13, 1) {real, imag} */,
  {32'hc5143ef8, 32'h00000000} /* (12, 13, 0) {real, imag} */,
  {32'hc52a58cd, 32'hc2617d50} /* (12, 12, 31) {real, imag} */,
  {32'h4485598e, 32'hc2bebf0a} /* (12, 12, 30) {real, imag} */,
  {32'hc24c0223, 32'h4229de97} /* (12, 12, 29) {real, imag} */,
  {32'hc24c5052, 32'h4372cc84} /* (12, 12, 28) {real, imag} */,
  {32'h4315a5de, 32'hc20e7e88} /* (12, 12, 27) {real, imag} */,
  {32'h42756748, 32'h41b6d3b1} /* (12, 12, 26) {real, imag} */,
  {32'hc0feab08, 32'hc2b89063} /* (12, 12, 25) {real, imag} */,
  {32'h427aa519, 32'hc1ce50da} /* (12, 12, 24) {real, imag} */,
  {32'h42a574a1, 32'h43067210} /* (12, 12, 23) {real, imag} */,
  {32'h4233282c, 32'h42c01637} /* (12, 12, 22) {real, imag} */,
  {32'hc04eb9e0, 32'hc26f9283} /* (12, 12, 21) {real, imag} */,
  {32'h417f5746, 32'hc1f0a341} /* (12, 12, 20) {real, imag} */,
  {32'hc16c1e6a, 32'hc069cb40} /* (12, 12, 19) {real, imag} */,
  {32'h4257e6d6, 32'hc23e93f1} /* (12, 12, 18) {real, imag} */,
  {32'h41b2eba1, 32'hc1acb0f4} /* (12, 12, 17) {real, imag} */,
  {32'h4285014a, 32'h00000000} /* (12, 12, 16) {real, imag} */,
  {32'h41b2eba1, 32'h41acb0f4} /* (12, 12, 15) {real, imag} */,
  {32'h4257e6d6, 32'h423e93f1} /* (12, 12, 14) {real, imag} */,
  {32'hc16c1e6a, 32'h4069cb40} /* (12, 12, 13) {real, imag} */,
  {32'h417f5746, 32'h41f0a341} /* (12, 12, 12) {real, imag} */,
  {32'hc04eb9e0, 32'h426f9283} /* (12, 12, 11) {real, imag} */,
  {32'h4233282c, 32'hc2c01637} /* (12, 12, 10) {real, imag} */,
  {32'h42a574a1, 32'hc3067210} /* (12, 12, 9) {real, imag} */,
  {32'h427aa519, 32'h41ce50da} /* (12, 12, 8) {real, imag} */,
  {32'hc0feab08, 32'h42b89063} /* (12, 12, 7) {real, imag} */,
  {32'h42756748, 32'hc1b6d3b1} /* (12, 12, 6) {real, imag} */,
  {32'h4315a5de, 32'h420e7e88} /* (12, 12, 5) {real, imag} */,
  {32'hc24c5052, 32'hc372cc84} /* (12, 12, 4) {real, imag} */,
  {32'hc24c0223, 32'hc229de97} /* (12, 12, 3) {real, imag} */,
  {32'h4485598e, 32'h42bebf0a} /* (12, 12, 2) {real, imag} */,
  {32'hc52a58cd, 32'h42617d50} /* (12, 12, 1) {real, imag} */,
  {32'hc4c60e37, 32'h00000000} /* (12, 12, 0) {real, imag} */,
  {32'hc4a7e048, 32'hc3bef370} /* (12, 11, 31) {real, imag} */,
  {32'h4427fb40, 32'hc2c6f88c} /* (12, 11, 30) {real, imag} */,
  {32'hc21c17c3, 32'h41e38241} /* (12, 11, 29) {real, imag} */,
  {32'hc3416198, 32'h42b93cde} /* (12, 11, 28) {real, imag} */,
  {32'h430f6d1a, 32'hc102b71c} /* (12, 11, 27) {real, imag} */,
  {32'hc267fd0c, 32'hc18d37f3} /* (12, 11, 26) {real, imag} */,
  {32'hc2e30d0e, 32'hc247b4b0} /* (12, 11, 25) {real, imag} */,
  {32'hc0d2f280, 32'hc1e50464} /* (12, 11, 24) {real, imag} */,
  {32'h42fef6da, 32'hc09eb7ca} /* (12, 11, 23) {real, imag} */,
  {32'h3ffd4278, 32'h41093528} /* (12, 11, 22) {real, imag} */,
  {32'hbe274f00, 32'hc30aed68} /* (12, 11, 21) {real, imag} */,
  {32'h42624eb4, 32'hc1c81030} /* (12, 11, 20) {real, imag} */,
  {32'h4183c1c8, 32'h3e9f3940} /* (12, 11, 19) {real, imag} */,
  {32'hc22b3280, 32'hc2600ab4} /* (12, 11, 18) {real, imag} */,
  {32'hc233e1e8, 32'hc1872caa} /* (12, 11, 17) {real, imag} */,
  {32'hc24ccb0a, 32'h00000000} /* (12, 11, 16) {real, imag} */,
  {32'hc233e1e8, 32'h41872caa} /* (12, 11, 15) {real, imag} */,
  {32'hc22b3280, 32'h42600ab4} /* (12, 11, 14) {real, imag} */,
  {32'h4183c1c8, 32'hbe9f3940} /* (12, 11, 13) {real, imag} */,
  {32'h42624eb4, 32'h41c81030} /* (12, 11, 12) {real, imag} */,
  {32'hbe274f00, 32'h430aed68} /* (12, 11, 11) {real, imag} */,
  {32'h3ffd4278, 32'hc1093528} /* (12, 11, 10) {real, imag} */,
  {32'h42fef6da, 32'h409eb7ca} /* (12, 11, 9) {real, imag} */,
  {32'hc0d2f280, 32'h41e50464} /* (12, 11, 8) {real, imag} */,
  {32'hc2e30d0e, 32'h4247b4b0} /* (12, 11, 7) {real, imag} */,
  {32'hc267fd0c, 32'h418d37f3} /* (12, 11, 6) {real, imag} */,
  {32'h430f6d1a, 32'h4102b71c} /* (12, 11, 5) {real, imag} */,
  {32'hc3416198, 32'hc2b93cde} /* (12, 11, 4) {real, imag} */,
  {32'hc21c17c3, 32'hc1e38241} /* (12, 11, 3) {real, imag} */,
  {32'h4427fb40, 32'h42c6f88c} /* (12, 11, 2) {real, imag} */,
  {32'hc4a7e048, 32'h43bef370} /* (12, 11, 1) {real, imag} */,
  {32'hc3bd3d1a, 32'h00000000} /* (12, 11, 0) {real, imag} */,
  {32'h44032b2f, 32'hc40d2dc0} /* (12, 10, 31) {real, imag} */,
  {32'hc2d05c28, 32'h4297e4b4} /* (12, 10, 30) {real, imag} */,
  {32'hc33d5562, 32'h412da794} /* (12, 10, 29) {real, imag} */,
  {32'hc20d48b8, 32'hc1ab1dc0} /* (12, 10, 28) {real, imag} */,
  {32'h42214f78, 32'h41d74180} /* (12, 10, 27) {real, imag} */,
  {32'h42298a38, 32'h4244ac49} /* (12, 10, 26) {real, imag} */,
  {32'h42c89c1b, 32'h4154282c} /* (12, 10, 25) {real, imag} */,
  {32'h4279be70, 32'h42940c50} /* (12, 10, 24) {real, imag} */,
  {32'hc1543080, 32'h41e38894} /* (12, 10, 23) {real, imag} */,
  {32'hc2fae425, 32'h420d0be0} /* (12, 10, 22) {real, imag} */,
  {32'hc2382064, 32'h3fcac050} /* (12, 10, 21) {real, imag} */,
  {32'h414ff688, 32'h42801dec} /* (12, 10, 20) {real, imag} */,
  {32'h42e095ff, 32'hc25b0884} /* (12, 10, 19) {real, imag} */,
  {32'h41b5426c, 32'h42d19595} /* (12, 10, 18) {real, imag} */,
  {32'hc1eb2067, 32'hc16ed289} /* (12, 10, 17) {real, imag} */,
  {32'hc12df750, 32'h00000000} /* (12, 10, 16) {real, imag} */,
  {32'hc1eb2067, 32'h416ed289} /* (12, 10, 15) {real, imag} */,
  {32'h41b5426c, 32'hc2d19595} /* (12, 10, 14) {real, imag} */,
  {32'h42e095ff, 32'h425b0884} /* (12, 10, 13) {real, imag} */,
  {32'h414ff688, 32'hc2801dec} /* (12, 10, 12) {real, imag} */,
  {32'hc2382064, 32'hbfcac050} /* (12, 10, 11) {real, imag} */,
  {32'hc2fae425, 32'hc20d0be0} /* (12, 10, 10) {real, imag} */,
  {32'hc1543080, 32'hc1e38894} /* (12, 10, 9) {real, imag} */,
  {32'h4279be70, 32'hc2940c50} /* (12, 10, 8) {real, imag} */,
  {32'h42c89c1b, 32'hc154282c} /* (12, 10, 7) {real, imag} */,
  {32'h42298a38, 32'hc244ac49} /* (12, 10, 6) {real, imag} */,
  {32'h42214f78, 32'hc1d74180} /* (12, 10, 5) {real, imag} */,
  {32'hc20d48b8, 32'h41ab1dc0} /* (12, 10, 4) {real, imag} */,
  {32'hc33d5562, 32'hc12da794} /* (12, 10, 3) {real, imag} */,
  {32'hc2d05c28, 32'hc297e4b4} /* (12, 10, 2) {real, imag} */,
  {32'h44032b2f, 32'h440d2dc0} /* (12, 10, 1) {real, imag} */,
  {32'h4494d5db, 32'h00000000} /* (12, 10, 0) {real, imag} */,
  {32'h44d7d9d2, 32'hc46ecea6} /* (12, 9, 31) {real, imag} */,
  {32'hc4458c21, 32'h437568fd} /* (12, 9, 30) {real, imag} */,
  {32'hc2a2aab1, 32'hc26516f6} /* (12, 9, 29) {real, imag} */,
  {32'h42d8df02, 32'hc1b0e5d8} /* (12, 9, 28) {real, imag} */,
  {32'hc251782c, 32'h42cf0d18} /* (12, 9, 27) {real, imag} */,
  {32'h416ff214, 32'h4113ddfe} /* (12, 9, 26) {real, imag} */,
  {32'h422856c4, 32'h41ab57e4} /* (12, 9, 25) {real, imag} */,
  {32'h41fab33d, 32'h42413d86} /* (12, 9, 24) {real, imag} */,
  {32'hc0fe01c8, 32'h3d9a3400} /* (12, 9, 23) {real, imag} */,
  {32'hc2a85936, 32'hc264d036} /* (12, 9, 22) {real, imag} */,
  {32'hc10f6e9c, 32'h40dca45c} /* (12, 9, 21) {real, imag} */,
  {32'hc20c97ac, 32'h3fe08340} /* (12, 9, 20) {real, imag} */,
  {32'hc1b43345, 32'h42638dea} /* (12, 9, 19) {real, imag} */,
  {32'hc29b33aa, 32'h42888ca6} /* (12, 9, 18) {real, imag} */,
  {32'hc1e7efa3, 32'h41766c7a} /* (12, 9, 17) {real, imag} */,
  {32'hc13a550b, 32'h00000000} /* (12, 9, 16) {real, imag} */,
  {32'hc1e7efa3, 32'hc1766c7a} /* (12, 9, 15) {real, imag} */,
  {32'hc29b33aa, 32'hc2888ca6} /* (12, 9, 14) {real, imag} */,
  {32'hc1b43345, 32'hc2638dea} /* (12, 9, 13) {real, imag} */,
  {32'hc20c97ac, 32'hbfe08340} /* (12, 9, 12) {real, imag} */,
  {32'hc10f6e9c, 32'hc0dca45c} /* (12, 9, 11) {real, imag} */,
  {32'hc2a85936, 32'h4264d036} /* (12, 9, 10) {real, imag} */,
  {32'hc0fe01c8, 32'hbd9a3400} /* (12, 9, 9) {real, imag} */,
  {32'h41fab33d, 32'hc2413d86} /* (12, 9, 8) {real, imag} */,
  {32'h422856c4, 32'hc1ab57e4} /* (12, 9, 7) {real, imag} */,
  {32'h416ff214, 32'hc113ddfe} /* (12, 9, 6) {real, imag} */,
  {32'hc251782c, 32'hc2cf0d18} /* (12, 9, 5) {real, imag} */,
  {32'h42d8df02, 32'h41b0e5d8} /* (12, 9, 4) {real, imag} */,
  {32'hc2a2aab1, 32'h426516f6} /* (12, 9, 3) {real, imag} */,
  {32'hc4458c21, 32'hc37568fd} /* (12, 9, 2) {real, imag} */,
  {32'h44d7d9d2, 32'h446ecea6} /* (12, 9, 1) {real, imag} */,
  {32'h450f6fc7, 32'h00000000} /* (12, 9, 0) {real, imag} */,
  {32'h4518b00e, 32'hc4a86951} /* (12, 8, 31) {real, imag} */,
  {32'hc48d1383, 32'h43b8aa0d} /* (12, 8, 30) {real, imag} */,
  {32'hc118c42c, 32'h400d02b0} /* (12, 8, 29) {real, imag} */,
  {32'h42921f54, 32'hc1803d20} /* (12, 8, 28) {real, imag} */,
  {32'hc28ca2ed, 32'hc15604d0} /* (12, 8, 27) {real, imag} */,
  {32'hc2088ffa, 32'h42995f14} /* (12, 8, 26) {real, imag} */,
  {32'h42ba8aa0, 32'hc16ef97a} /* (12, 8, 25) {real, imag} */,
  {32'h42851e5c, 32'h426bb588} /* (12, 8, 24) {real, imag} */,
  {32'h414b591c, 32'hc2da00a7} /* (12, 8, 23) {real, imag} */,
  {32'hc1b171f8, 32'h4252e765} /* (12, 8, 22) {real, imag} */,
  {32'hc21eaa25, 32'h42c227f7} /* (12, 8, 21) {real, imag} */,
  {32'h42ab1ff1, 32'hc2b99c77} /* (12, 8, 20) {real, imag} */,
  {32'hc30df228, 32'hc282181b} /* (12, 8, 19) {real, imag} */,
  {32'hc235d4e2, 32'h43006396} /* (12, 8, 18) {real, imag} */,
  {32'h41e2c23d, 32'h4231466a} /* (12, 8, 17) {real, imag} */,
  {32'h42258655, 32'h00000000} /* (12, 8, 16) {real, imag} */,
  {32'h41e2c23d, 32'hc231466a} /* (12, 8, 15) {real, imag} */,
  {32'hc235d4e2, 32'hc3006396} /* (12, 8, 14) {real, imag} */,
  {32'hc30df228, 32'h4282181b} /* (12, 8, 13) {real, imag} */,
  {32'h42ab1ff1, 32'h42b99c77} /* (12, 8, 12) {real, imag} */,
  {32'hc21eaa25, 32'hc2c227f7} /* (12, 8, 11) {real, imag} */,
  {32'hc1b171f8, 32'hc252e765} /* (12, 8, 10) {real, imag} */,
  {32'h414b591c, 32'h42da00a7} /* (12, 8, 9) {real, imag} */,
  {32'h42851e5c, 32'hc26bb588} /* (12, 8, 8) {real, imag} */,
  {32'h42ba8aa0, 32'h416ef97a} /* (12, 8, 7) {real, imag} */,
  {32'hc2088ffa, 32'hc2995f14} /* (12, 8, 6) {real, imag} */,
  {32'hc28ca2ed, 32'h415604d0} /* (12, 8, 5) {real, imag} */,
  {32'h42921f54, 32'h41803d20} /* (12, 8, 4) {real, imag} */,
  {32'hc118c42c, 32'hc00d02b0} /* (12, 8, 3) {real, imag} */,
  {32'hc48d1383, 32'hc3b8aa0d} /* (12, 8, 2) {real, imag} */,
  {32'h4518b00e, 32'h44a86951} /* (12, 8, 1) {real, imag} */,
  {32'h45459d50, 32'h00000000} /* (12, 8, 0) {real, imag} */,
  {32'h453e2617, 32'hc4c2854b} /* (12, 7, 31) {real, imag} */,
  {32'hc480ffb2, 32'h442e5b4e} /* (12, 7, 30) {real, imag} */,
  {32'hc266e1be, 32'h4199dce3} /* (12, 7, 29) {real, imag} */,
  {32'h4225e830, 32'hc1cb8c36} /* (12, 7, 28) {real, imag} */,
  {32'hc34efa0d, 32'h42e42cd6} /* (12, 7, 27) {real, imag} */,
  {32'hc1379c70, 32'hc0d60020} /* (12, 7, 26) {real, imag} */,
  {32'h4279df14, 32'hc318d811} /* (12, 7, 25) {real, imag} */,
  {32'hc14ba194, 32'h42f23279} /* (12, 7, 24) {real, imag} */,
  {32'h42712840, 32'hc2846928} /* (12, 7, 23) {real, imag} */,
  {32'hc21e3680, 32'h4338246d} /* (12, 7, 22) {real, imag} */,
  {32'hc2fa98d2, 32'h423cd110} /* (12, 7, 21) {real, imag} */,
  {32'h42098933, 32'h4026bc60} /* (12, 7, 20) {real, imag} */,
  {32'hc233649f, 32'h41c61e58} /* (12, 7, 19) {real, imag} */,
  {32'hc227531e, 32'hc1ea7c4b} /* (12, 7, 18) {real, imag} */,
  {32'h41b3dd4c, 32'hc2bfcdec} /* (12, 7, 17) {real, imag} */,
  {32'h429d9584, 32'h00000000} /* (12, 7, 16) {real, imag} */,
  {32'h41b3dd4c, 32'h42bfcdec} /* (12, 7, 15) {real, imag} */,
  {32'hc227531e, 32'h41ea7c4b} /* (12, 7, 14) {real, imag} */,
  {32'hc233649f, 32'hc1c61e58} /* (12, 7, 13) {real, imag} */,
  {32'h42098933, 32'hc026bc60} /* (12, 7, 12) {real, imag} */,
  {32'hc2fa98d2, 32'hc23cd110} /* (12, 7, 11) {real, imag} */,
  {32'hc21e3680, 32'hc338246d} /* (12, 7, 10) {real, imag} */,
  {32'h42712840, 32'h42846928} /* (12, 7, 9) {real, imag} */,
  {32'hc14ba194, 32'hc2f23279} /* (12, 7, 8) {real, imag} */,
  {32'h4279df14, 32'h4318d811} /* (12, 7, 7) {real, imag} */,
  {32'hc1379c70, 32'h40d60020} /* (12, 7, 6) {real, imag} */,
  {32'hc34efa0d, 32'hc2e42cd6} /* (12, 7, 5) {real, imag} */,
  {32'h4225e830, 32'h41cb8c36} /* (12, 7, 4) {real, imag} */,
  {32'hc266e1be, 32'hc199dce3} /* (12, 7, 3) {real, imag} */,
  {32'hc480ffb2, 32'hc42e5b4e} /* (12, 7, 2) {real, imag} */,
  {32'h453e2617, 32'h44c2854b} /* (12, 7, 1) {real, imag} */,
  {32'h456419cd, 32'h00000000} /* (12, 7, 0) {real, imag} */,
  {32'h454822df, 32'hc503120f} /* (12, 6, 31) {real, imag} */,
  {32'hc456e734, 32'h446156a6} /* (12, 6, 30) {real, imag} */,
  {32'hc2527f4a, 32'h42911164} /* (12, 6, 29) {real, imag} */,
  {32'h41f5dc50, 32'h423a2e6c} /* (12, 6, 28) {real, imag} */,
  {32'hc2bfccbc, 32'h435d57c3} /* (12, 6, 27) {real, imag} */,
  {32'hc206d749, 32'h41ce791a} /* (12, 6, 26) {real, imag} */,
  {32'hc28471e3, 32'hc29a7386} /* (12, 6, 25) {real, imag} */,
  {32'hc19687c1, 32'h41bc665c} /* (12, 6, 24) {real, imag} */,
  {32'h421d540c, 32'h42b189b4} /* (12, 6, 23) {real, imag} */,
  {32'hc2af6567, 32'hc28edd93} /* (12, 6, 22) {real, imag} */,
  {32'h41a4ecc6, 32'hc104cc90} /* (12, 6, 21) {real, imag} */,
  {32'hc22fcd4f, 32'hc241136e} /* (12, 6, 20) {real, imag} */,
  {32'h4280840c, 32'h41de3afe} /* (12, 6, 19) {real, imag} */,
  {32'hc2bdab36, 32'h4176e524} /* (12, 6, 18) {real, imag} */,
  {32'h42815cce, 32'hc083f24a} /* (12, 6, 17) {real, imag} */,
  {32'hc2ab2299, 32'h00000000} /* (12, 6, 16) {real, imag} */,
  {32'h42815cce, 32'h4083f24a} /* (12, 6, 15) {real, imag} */,
  {32'hc2bdab36, 32'hc176e524} /* (12, 6, 14) {real, imag} */,
  {32'h4280840c, 32'hc1de3afe} /* (12, 6, 13) {real, imag} */,
  {32'hc22fcd4f, 32'h4241136e} /* (12, 6, 12) {real, imag} */,
  {32'h41a4ecc6, 32'h4104cc90} /* (12, 6, 11) {real, imag} */,
  {32'hc2af6567, 32'h428edd93} /* (12, 6, 10) {real, imag} */,
  {32'h421d540c, 32'hc2b189b4} /* (12, 6, 9) {real, imag} */,
  {32'hc19687c1, 32'hc1bc665c} /* (12, 6, 8) {real, imag} */,
  {32'hc28471e3, 32'h429a7386} /* (12, 6, 7) {real, imag} */,
  {32'hc206d749, 32'hc1ce791a} /* (12, 6, 6) {real, imag} */,
  {32'hc2bfccbc, 32'hc35d57c3} /* (12, 6, 5) {real, imag} */,
  {32'h41f5dc50, 32'hc23a2e6c} /* (12, 6, 4) {real, imag} */,
  {32'hc2527f4a, 32'hc2911164} /* (12, 6, 3) {real, imag} */,
  {32'hc456e734, 32'hc46156a6} /* (12, 6, 2) {real, imag} */,
  {32'h454822df, 32'h4503120f} /* (12, 6, 1) {real, imag} */,
  {32'h4581e0b4, 32'h00000000} /* (12, 6, 0) {real, imag} */,
  {32'h453cc780, 32'hc5344f84} /* (12, 5, 31) {real, imag} */,
  {32'hc398da8c, 32'h44768e20} /* (12, 5, 30) {real, imag} */,
  {32'hc31bc4dc, 32'h419560a9} /* (12, 5, 29) {real, imag} */,
  {32'hc232d10e, 32'h43307685} /* (12, 5, 28) {real, imag} */,
  {32'hc3344a30, 32'h42267845} /* (12, 5, 27) {real, imag} */,
  {32'hc2b6fd54, 32'h42e42a66} /* (12, 5, 26) {real, imag} */,
  {32'h4246b376, 32'hc258d756} /* (12, 5, 25) {real, imag} */,
  {32'h402da780, 32'h42c4dcf5} /* (12, 5, 24) {real, imag} */,
  {32'hc1e36bea, 32'hc2aa9f78} /* (12, 5, 23) {real, imag} */,
  {32'h40d8fad6, 32'h42691ae2} /* (12, 5, 22) {real, imag} */,
  {32'h426da40d, 32'hc2214106} /* (12, 5, 21) {real, imag} */,
  {32'hc1347390, 32'hc239b718} /* (12, 5, 20) {real, imag} */,
  {32'hc07be420, 32'h424ad4f2} /* (12, 5, 19) {real, imag} */,
  {32'h410d7542, 32'h423cb2d8} /* (12, 5, 18) {real, imag} */,
  {32'hc2057f76, 32'hc267ecd4} /* (12, 5, 17) {real, imag} */,
  {32'hc102c3a6, 32'h00000000} /* (12, 5, 16) {real, imag} */,
  {32'hc2057f76, 32'h4267ecd4} /* (12, 5, 15) {real, imag} */,
  {32'h410d7542, 32'hc23cb2d8} /* (12, 5, 14) {real, imag} */,
  {32'hc07be420, 32'hc24ad4f2} /* (12, 5, 13) {real, imag} */,
  {32'hc1347390, 32'h4239b718} /* (12, 5, 12) {real, imag} */,
  {32'h426da40d, 32'h42214106} /* (12, 5, 11) {real, imag} */,
  {32'h40d8fad6, 32'hc2691ae2} /* (12, 5, 10) {real, imag} */,
  {32'hc1e36bea, 32'h42aa9f78} /* (12, 5, 9) {real, imag} */,
  {32'h402da780, 32'hc2c4dcf5} /* (12, 5, 8) {real, imag} */,
  {32'h4246b376, 32'h4258d756} /* (12, 5, 7) {real, imag} */,
  {32'hc2b6fd54, 32'hc2e42a66} /* (12, 5, 6) {real, imag} */,
  {32'hc3344a30, 32'hc2267845} /* (12, 5, 5) {real, imag} */,
  {32'hc232d10e, 32'hc3307685} /* (12, 5, 4) {real, imag} */,
  {32'hc31bc4dc, 32'hc19560a9} /* (12, 5, 3) {real, imag} */,
  {32'hc398da8c, 32'hc4768e20} /* (12, 5, 2) {real, imag} */,
  {32'h453cc780, 32'h45344f84} /* (12, 5, 1) {real, imag} */,
  {32'h459475cf, 32'h00000000} /* (12, 5, 0) {real, imag} */,
  {32'h45329f66, 32'hc55a9417} /* (12, 4, 31) {real, imag} */,
  {32'h42c0d148, 32'h448d91c8} /* (12, 4, 30) {real, imag} */,
  {32'hc2dec352, 32'hc25a6067} /* (12, 4, 29) {real, imag} */,
  {32'hc319733e, 32'h435dbe73} /* (12, 4, 28) {real, imag} */,
  {32'hc321f723, 32'hc095957a} /* (12, 4, 27) {real, imag} */,
  {32'hc04b2ecc, 32'h4250de60} /* (12, 4, 26) {real, imag} */,
  {32'hc27c11d5, 32'hc3115aac} /* (12, 4, 25) {real, imag} */,
  {32'hc22dc94e, 32'h4284047f} /* (12, 4, 24) {real, imag} */,
  {32'hc2118c63, 32'h42297ae8} /* (12, 4, 23) {real, imag} */,
  {32'hc298e930, 32'h42bc38be} /* (12, 4, 22) {real, imag} */,
  {32'h41a33f13, 32'h428a50e2} /* (12, 4, 21) {real, imag} */,
  {32'hc163042d, 32'hc03e72d8} /* (12, 4, 20) {real, imag} */,
  {32'hc1e2a060, 32'h42302edc} /* (12, 4, 19) {real, imag} */,
  {32'h42a34903, 32'hc27f3678} /* (12, 4, 18) {real, imag} */,
  {32'hc0e91748, 32'hc22888fc} /* (12, 4, 17) {real, imag} */,
  {32'hc161e553, 32'h00000000} /* (12, 4, 16) {real, imag} */,
  {32'hc0e91748, 32'h422888fc} /* (12, 4, 15) {real, imag} */,
  {32'h42a34903, 32'h427f3678} /* (12, 4, 14) {real, imag} */,
  {32'hc1e2a060, 32'hc2302edc} /* (12, 4, 13) {real, imag} */,
  {32'hc163042d, 32'h403e72d8} /* (12, 4, 12) {real, imag} */,
  {32'h41a33f13, 32'hc28a50e2} /* (12, 4, 11) {real, imag} */,
  {32'hc298e930, 32'hc2bc38be} /* (12, 4, 10) {real, imag} */,
  {32'hc2118c63, 32'hc2297ae8} /* (12, 4, 9) {real, imag} */,
  {32'hc22dc94e, 32'hc284047f} /* (12, 4, 8) {real, imag} */,
  {32'hc27c11d5, 32'h43115aac} /* (12, 4, 7) {real, imag} */,
  {32'hc04b2ecc, 32'hc250de60} /* (12, 4, 6) {real, imag} */,
  {32'hc321f723, 32'h4095957a} /* (12, 4, 5) {real, imag} */,
  {32'hc319733e, 32'hc35dbe73} /* (12, 4, 4) {real, imag} */,
  {32'hc2dec352, 32'h425a6067} /* (12, 4, 3) {real, imag} */,
  {32'h42c0d148, 32'hc48d91c8} /* (12, 4, 2) {real, imag} */,
  {32'h45329f66, 32'h455a9417} /* (12, 4, 1) {real, imag} */,
  {32'h459d5885, 32'h00000000} /* (12, 4, 0) {real, imag} */,
  {32'h452f6746, 32'hc566e0d6} /* (12, 3, 31) {real, imag} */,
  {32'h43584dd8, 32'h448a072c} /* (12, 3, 30) {real, imag} */,
  {32'hc2439e5e, 32'h4286a304} /* (12, 3, 29) {real, imag} */,
  {32'hc350dcae, 32'h42d2ac4a} /* (12, 3, 28) {real, imag} */,
  {32'hc38caebd, 32'hc33b0c58} /* (12, 3, 27) {real, imag} */,
  {32'hc29efbe4, 32'h4219fb18} /* (12, 3, 26) {real, imag} */,
  {32'h4150414c, 32'hc2c540d6} /* (12, 3, 25) {real, imag} */,
  {32'h4236975d, 32'h431fdb4d} /* (12, 3, 24) {real, imag} */,
  {32'hc1d7fd9a, 32'h42f32f41} /* (12, 3, 23) {real, imag} */,
  {32'hc0d84ef0, 32'h42b2fc14} /* (12, 3, 22) {real, imag} */,
  {32'hc30f8c18, 32'hc1e4a8bd} /* (12, 3, 21) {real, imag} */,
  {32'hc030c850, 32'hc28ebb6d} /* (12, 3, 20) {real, imag} */,
  {32'h42490af7, 32'hc286a1a0} /* (12, 3, 19) {real, imag} */,
  {32'h425c1843, 32'hc2980de6} /* (12, 3, 18) {real, imag} */,
  {32'hc1b1ec21, 32'h421d3450} /* (12, 3, 17) {real, imag} */,
  {32'hc236538e, 32'h00000000} /* (12, 3, 16) {real, imag} */,
  {32'hc1b1ec21, 32'hc21d3450} /* (12, 3, 15) {real, imag} */,
  {32'h425c1843, 32'h42980de6} /* (12, 3, 14) {real, imag} */,
  {32'h42490af7, 32'h4286a1a0} /* (12, 3, 13) {real, imag} */,
  {32'hc030c850, 32'h428ebb6d} /* (12, 3, 12) {real, imag} */,
  {32'hc30f8c18, 32'h41e4a8bd} /* (12, 3, 11) {real, imag} */,
  {32'hc0d84ef0, 32'hc2b2fc14} /* (12, 3, 10) {real, imag} */,
  {32'hc1d7fd9a, 32'hc2f32f41} /* (12, 3, 9) {real, imag} */,
  {32'h4236975d, 32'hc31fdb4d} /* (12, 3, 8) {real, imag} */,
  {32'h4150414c, 32'h42c540d6} /* (12, 3, 7) {real, imag} */,
  {32'hc29efbe4, 32'hc219fb18} /* (12, 3, 6) {real, imag} */,
  {32'hc38caebd, 32'h433b0c58} /* (12, 3, 5) {real, imag} */,
  {32'hc350dcae, 32'hc2d2ac4a} /* (12, 3, 4) {real, imag} */,
  {32'hc2439e5e, 32'hc286a304} /* (12, 3, 3) {real, imag} */,
  {32'h43584dd8, 32'hc48a072c} /* (12, 3, 2) {real, imag} */,
  {32'h452f6746, 32'h4566e0d6} /* (12, 3, 1) {real, imag} */,
  {32'h459ee0f3, 32'h00000000} /* (12, 3, 0) {real, imag} */,
  {32'h453760de, 32'hc56741bf} /* (12, 2, 31) {real, imag} */,
  {32'h434fef2c, 32'h4484beb1} /* (12, 2, 30) {real, imag} */,
  {32'hc3379a89, 32'h430e763e} /* (12, 2, 29) {real, imag} */,
  {32'hc20d36ed, 32'h438c8b66} /* (12, 2, 28) {real, imag} */,
  {32'hc36113e8, 32'hc35815d4} /* (12, 2, 27) {real, imag} */,
  {32'hc2bd77de, 32'hc2d44e3b} /* (12, 2, 26) {real, imag} */,
  {32'h428b27a3, 32'h43010385} /* (12, 2, 25) {real, imag} */,
  {32'h42c90ff5, 32'hc1dcc79a} /* (12, 2, 24) {real, imag} */,
  {32'h40271e28, 32'h427bc4a0} /* (12, 2, 23) {real, imag} */,
  {32'hc1b0fd5b, 32'h4270cbb2} /* (12, 2, 22) {real, imag} */,
  {32'hc2d1abe5, 32'hc06fe4fc} /* (12, 2, 21) {real, imag} */,
  {32'hc30ccea4, 32'h421e61ae} /* (12, 2, 20) {real, imag} */,
  {32'hc1f1303d, 32'h41b5f6ca} /* (12, 2, 19) {real, imag} */,
  {32'h42cba75d, 32'hc2bde6c2} /* (12, 2, 18) {real, imag} */,
  {32'hc269e379, 32'h4139cea8} /* (12, 2, 17) {real, imag} */,
  {32'h4232a3a9, 32'h00000000} /* (12, 2, 16) {real, imag} */,
  {32'hc269e379, 32'hc139cea8} /* (12, 2, 15) {real, imag} */,
  {32'h42cba75d, 32'h42bde6c2} /* (12, 2, 14) {real, imag} */,
  {32'hc1f1303d, 32'hc1b5f6ca} /* (12, 2, 13) {real, imag} */,
  {32'hc30ccea4, 32'hc21e61ae} /* (12, 2, 12) {real, imag} */,
  {32'hc2d1abe5, 32'h406fe4fc} /* (12, 2, 11) {real, imag} */,
  {32'hc1b0fd5b, 32'hc270cbb2} /* (12, 2, 10) {real, imag} */,
  {32'h40271e28, 32'hc27bc4a0} /* (12, 2, 9) {real, imag} */,
  {32'h42c90ff5, 32'h41dcc79a} /* (12, 2, 8) {real, imag} */,
  {32'h428b27a3, 32'hc3010385} /* (12, 2, 7) {real, imag} */,
  {32'hc2bd77de, 32'h42d44e3b} /* (12, 2, 6) {real, imag} */,
  {32'hc36113e8, 32'h435815d4} /* (12, 2, 5) {real, imag} */,
  {32'hc20d36ed, 32'hc38c8b66} /* (12, 2, 4) {real, imag} */,
  {32'hc3379a89, 32'hc30e763e} /* (12, 2, 3) {real, imag} */,
  {32'h434fef2c, 32'hc484beb1} /* (12, 2, 2) {real, imag} */,
  {32'h453760de, 32'h456741bf} /* (12, 2, 1) {real, imag} */,
  {32'h45a3092f, 32'h00000000} /* (12, 2, 0) {real, imag} */,
  {32'h453d4878, 32'hc557b7e6} /* (12, 1, 31) {real, imag} */,
  {32'h42e6732c, 32'h4475a3bc} /* (12, 1, 30) {real, imag} */,
  {32'hc13b2f38, 32'h4218c204} /* (12, 1, 29) {real, imag} */,
  {32'hc2476dc5, 32'h43c6b49a} /* (12, 1, 28) {real, imag} */,
  {32'hc30f828a, 32'hc37f90f6} /* (12, 1, 27) {real, imag} */,
  {32'h4237e3ba, 32'hc1d1d58e} /* (12, 1, 26) {real, imag} */,
  {32'hc0b1f5c8, 32'h3fab81e8} /* (12, 1, 25) {real, imag} */,
  {32'h42f7f591, 32'hc108c313} /* (12, 1, 24) {real, imag} */,
  {32'hc25469b2, 32'hc0e49f48} /* (12, 1, 23) {real, imag} */,
  {32'hc275e322, 32'h42a79224} /* (12, 1, 22) {real, imag} */,
  {32'h40af02a8, 32'h42bfee74} /* (12, 1, 21) {real, imag} */,
  {32'hc156c224, 32'hbff747b0} /* (12, 1, 20) {real, imag} */,
  {32'hc29c3c93, 32'h428c57bb} /* (12, 1, 19) {real, imag} */,
  {32'h424923a0, 32'hc2a0767f} /* (12, 1, 18) {real, imag} */,
  {32'hc2028754, 32'h41a865fa} /* (12, 1, 17) {real, imag} */,
  {32'hc18133cf, 32'h00000000} /* (12, 1, 16) {real, imag} */,
  {32'hc2028754, 32'hc1a865fa} /* (12, 1, 15) {real, imag} */,
  {32'h424923a0, 32'h42a0767f} /* (12, 1, 14) {real, imag} */,
  {32'hc29c3c93, 32'hc28c57bb} /* (12, 1, 13) {real, imag} */,
  {32'hc156c224, 32'h3ff747b0} /* (12, 1, 12) {real, imag} */,
  {32'h40af02a8, 32'hc2bfee74} /* (12, 1, 11) {real, imag} */,
  {32'hc275e322, 32'hc2a79224} /* (12, 1, 10) {real, imag} */,
  {32'hc25469b2, 32'h40e49f48} /* (12, 1, 9) {real, imag} */,
  {32'h42f7f591, 32'h4108c313} /* (12, 1, 8) {real, imag} */,
  {32'hc0b1f5c8, 32'hbfab81e8} /* (12, 1, 7) {real, imag} */,
  {32'h4237e3ba, 32'h41d1d58e} /* (12, 1, 6) {real, imag} */,
  {32'hc30f828a, 32'h437f90f6} /* (12, 1, 5) {real, imag} */,
  {32'hc2476dc5, 32'hc3c6b49a} /* (12, 1, 4) {real, imag} */,
  {32'hc13b2f38, 32'hc218c204} /* (12, 1, 3) {real, imag} */,
  {32'h42e6732c, 32'hc475a3bc} /* (12, 1, 2) {real, imag} */,
  {32'h453d4878, 32'h4557b7e6} /* (12, 1, 1) {real, imag} */,
  {32'h459d5512, 32'h00000000} /* (12, 1, 0) {real, imag} */,
  {32'h4544c76b, 32'hc52e1f7a} /* (12, 0, 31) {real, imag} */,
  {32'hc3a5ab4a, 32'h444609da} /* (12, 0, 30) {real, imag} */,
  {32'hc203fe81, 32'h41a4037a} /* (12, 0, 29) {real, imag} */,
  {32'hc29fe4ec, 32'h431d9537} /* (12, 0, 28) {real, imag} */,
  {32'hc309acfd, 32'hc304e283} /* (12, 0, 27) {real, imag} */,
  {32'hc158c004, 32'h41281081} /* (12, 0, 26) {real, imag} */,
  {32'h41916512, 32'hc2a1d93e} /* (12, 0, 25) {real, imag} */,
  {32'h428fa6ad, 32'hc1ae1f61} /* (12, 0, 24) {real, imag} */,
  {32'hc26d54e8, 32'h412d4df6} /* (12, 0, 23) {real, imag} */,
  {32'h4236a2e5, 32'h41cf0dda} /* (12, 0, 22) {real, imag} */,
  {32'h41bcdddd, 32'h40c86938} /* (12, 0, 21) {real, imag} */,
  {32'h41f72efe, 32'hc1de3644} /* (12, 0, 20) {real, imag} */,
  {32'hc129f64a, 32'h42874d10} /* (12, 0, 19) {real, imag} */,
  {32'h41a75f9e, 32'h420ba462} /* (12, 0, 18) {real, imag} */,
  {32'h422c2264, 32'h41bc1e9f} /* (12, 0, 17) {real, imag} */,
  {32'hc243449d, 32'h00000000} /* (12, 0, 16) {real, imag} */,
  {32'h422c2264, 32'hc1bc1e9f} /* (12, 0, 15) {real, imag} */,
  {32'h41a75f9e, 32'hc20ba462} /* (12, 0, 14) {real, imag} */,
  {32'hc129f64a, 32'hc2874d10} /* (12, 0, 13) {real, imag} */,
  {32'h41f72efe, 32'h41de3644} /* (12, 0, 12) {real, imag} */,
  {32'h41bcdddd, 32'hc0c86938} /* (12, 0, 11) {real, imag} */,
  {32'h4236a2e5, 32'hc1cf0dda} /* (12, 0, 10) {real, imag} */,
  {32'hc26d54e8, 32'hc12d4df6} /* (12, 0, 9) {real, imag} */,
  {32'h428fa6ad, 32'h41ae1f61} /* (12, 0, 8) {real, imag} */,
  {32'h41916512, 32'h42a1d93e} /* (12, 0, 7) {real, imag} */,
  {32'hc158c004, 32'hc1281081} /* (12, 0, 6) {real, imag} */,
  {32'hc309acfd, 32'h4304e283} /* (12, 0, 5) {real, imag} */,
  {32'hc29fe4ec, 32'hc31d9537} /* (12, 0, 4) {real, imag} */,
  {32'hc203fe81, 32'hc1a4037a} /* (12, 0, 3) {real, imag} */,
  {32'hc3a5ab4a, 32'hc44609da} /* (12, 0, 2) {real, imag} */,
  {32'h4544c76b, 32'h452e1f7a} /* (12, 0, 1) {real, imag} */,
  {32'h45984ff7, 32'h00000000} /* (12, 0, 0) {real, imag} */,
  {32'h4580b08d, 32'hc51085c2} /* (11, 31, 31) {real, imag} */,
  {32'hc456c99d, 32'h44379a39} /* (11, 31, 30) {real, imag} */,
  {32'hc2304cb4, 32'h421dedc0} /* (11, 31, 29) {real, imag} */,
  {32'h42957d51, 32'h42a3c13a} /* (11, 31, 28) {real, imag} */,
  {32'hc30bf696, 32'h41e7b6b0} /* (11, 31, 27) {real, imag} */,
  {32'hc19aee78, 32'hc1dabf22} /* (11, 31, 26) {real, imag} */,
  {32'h42ccc25e, 32'hc25f191c} /* (11, 31, 25) {real, imag} */,
  {32'hc2d4801f, 32'h4267c1e0} /* (11, 31, 24) {real, imag} */,
  {32'h3fe4da80, 32'hc207e114} /* (11, 31, 23) {real, imag} */,
  {32'h42054503, 32'h413e8d5c} /* (11, 31, 22) {real, imag} */,
  {32'h422054be, 32'h41999196} /* (11, 31, 21) {real, imag} */,
  {32'h41ded65b, 32'hc24c16ea} /* (11, 31, 20) {real, imag} */,
  {32'h42d2a29c, 32'hc2887d0f} /* (11, 31, 19) {real, imag} */,
  {32'h42232323, 32'h425aea96} /* (11, 31, 18) {real, imag} */,
  {32'h41b9c876, 32'hc2b0934e} /* (11, 31, 17) {real, imag} */,
  {32'h4309728f, 32'h00000000} /* (11, 31, 16) {real, imag} */,
  {32'h41b9c876, 32'h42b0934e} /* (11, 31, 15) {real, imag} */,
  {32'h42232323, 32'hc25aea96} /* (11, 31, 14) {real, imag} */,
  {32'h42d2a29c, 32'h42887d0f} /* (11, 31, 13) {real, imag} */,
  {32'h41ded65b, 32'h424c16ea} /* (11, 31, 12) {real, imag} */,
  {32'h422054be, 32'hc1999196} /* (11, 31, 11) {real, imag} */,
  {32'h42054503, 32'hc13e8d5c} /* (11, 31, 10) {real, imag} */,
  {32'h3fe4da80, 32'h4207e114} /* (11, 31, 9) {real, imag} */,
  {32'hc2d4801f, 32'hc267c1e0} /* (11, 31, 8) {real, imag} */,
  {32'h42ccc25e, 32'h425f191c} /* (11, 31, 7) {real, imag} */,
  {32'hc19aee78, 32'h41dabf22} /* (11, 31, 6) {real, imag} */,
  {32'hc30bf696, 32'hc1e7b6b0} /* (11, 31, 5) {real, imag} */,
  {32'h42957d51, 32'hc2a3c13a} /* (11, 31, 4) {real, imag} */,
  {32'hc2304cb4, 32'hc21dedc0} /* (11, 31, 3) {real, imag} */,
  {32'hc456c99d, 32'hc4379a39} /* (11, 31, 2) {real, imag} */,
  {32'h4580b08d, 32'h451085c2} /* (11, 31, 1) {real, imag} */,
  {32'h45a9f1cd, 32'h00000000} /* (11, 31, 0) {real, imag} */,
  {32'h458feef9, 32'hc4d98c4c} /* (11, 30, 31) {real, imag} */,
  {32'hc4ad3eae, 32'h44310ca8} /* (11, 30, 30) {real, imag} */,
  {32'hc1f26293, 32'h42ad15b2} /* (11, 30, 29) {real, imag} */,
  {32'h4297e14b, 32'h42a9ce3a} /* (11, 30, 28) {real, imag} */,
  {32'hc31f48e0, 32'hc2ab3c99} /* (11, 30, 27) {real, imag} */,
  {32'h41b0d48c, 32'hc31b1c58} /* (11, 30, 26) {real, imag} */,
  {32'h42608967, 32'h424c865b} /* (11, 30, 25) {real, imag} */,
  {32'hc1a9e22c, 32'hbfeca420} /* (11, 30, 24) {real, imag} */,
  {32'hc221224d, 32'hc2b9a630} /* (11, 30, 23) {real, imag} */,
  {32'h4213b73d, 32'hc1a4a33c} /* (11, 30, 22) {real, imag} */,
  {32'hc2b819de, 32'h4282f6e6} /* (11, 30, 21) {real, imag} */,
  {32'hc1d5efe8, 32'hc3035f9e} /* (11, 30, 20) {real, imag} */,
  {32'hc17847d0, 32'hc21a932f} /* (11, 30, 19) {real, imag} */,
  {32'h418a477a, 32'hc0a6c69a} /* (11, 30, 18) {real, imag} */,
  {32'h419144ad, 32'hc1826e21} /* (11, 30, 17) {real, imag} */,
  {32'h425edeb6, 32'h00000000} /* (11, 30, 16) {real, imag} */,
  {32'h419144ad, 32'h41826e21} /* (11, 30, 15) {real, imag} */,
  {32'h418a477a, 32'h40a6c69a} /* (11, 30, 14) {real, imag} */,
  {32'hc17847d0, 32'h421a932f} /* (11, 30, 13) {real, imag} */,
  {32'hc1d5efe8, 32'h43035f9e} /* (11, 30, 12) {real, imag} */,
  {32'hc2b819de, 32'hc282f6e6} /* (11, 30, 11) {real, imag} */,
  {32'h4213b73d, 32'h41a4a33c} /* (11, 30, 10) {real, imag} */,
  {32'hc221224d, 32'h42b9a630} /* (11, 30, 9) {real, imag} */,
  {32'hc1a9e22c, 32'h3feca420} /* (11, 30, 8) {real, imag} */,
  {32'h42608967, 32'hc24c865b} /* (11, 30, 7) {real, imag} */,
  {32'h41b0d48c, 32'h431b1c58} /* (11, 30, 6) {real, imag} */,
  {32'hc31f48e0, 32'h42ab3c99} /* (11, 30, 5) {real, imag} */,
  {32'h4297e14b, 32'hc2a9ce3a} /* (11, 30, 4) {real, imag} */,
  {32'hc1f26293, 32'hc2ad15b2} /* (11, 30, 3) {real, imag} */,
  {32'hc4ad3eae, 32'hc4310ca8} /* (11, 30, 2) {real, imag} */,
  {32'h458feef9, 32'h44d98c4c} /* (11, 30, 1) {real, imag} */,
  {32'h45b00b9b, 32'h00000000} /* (11, 30, 0) {real, imag} */,
  {32'h459892e6, 32'hc4b245c2} /* (11, 29, 31) {real, imag} */,
  {32'hc4b8fc2c, 32'h4408e4b9} /* (11, 29, 30) {real, imag} */,
  {32'h4233475d, 32'h3fab3c50} /* (11, 29, 29) {real, imag} */,
  {32'h43373972, 32'hc29b6327} /* (11, 29, 28) {real, imag} */,
  {32'hc3784552, 32'hc1e64ce9} /* (11, 29, 27) {real, imag} */,
  {32'h418a0b14, 32'hc24bacec} /* (11, 29, 26) {real, imag} */,
  {32'hc158b272, 32'h427a85f4} /* (11, 29, 25) {real, imag} */,
  {32'hc1ffffce, 32'h41dd7e6c} /* (11, 29, 24) {real, imag} */,
  {32'hc1d7de8c, 32'hc17b9dc4} /* (11, 29, 23) {real, imag} */,
  {32'h42465da2, 32'h41edbe04} /* (11, 29, 22) {real, imag} */,
  {32'hc206a812, 32'hc195ad96} /* (11, 29, 21) {real, imag} */,
  {32'hc125b563, 32'h41aa4e6a} /* (11, 29, 20) {real, imag} */,
  {32'hc27d4eae, 32'h4231b2c2} /* (11, 29, 19) {real, imag} */,
  {32'hc220c1c1, 32'h3fde2240} /* (11, 29, 18) {real, imag} */,
  {32'h41892ce4, 32'h4110533c} /* (11, 29, 17) {real, imag} */,
  {32'h42179d6e, 32'h00000000} /* (11, 29, 16) {real, imag} */,
  {32'h41892ce4, 32'hc110533c} /* (11, 29, 15) {real, imag} */,
  {32'hc220c1c1, 32'hbfde2240} /* (11, 29, 14) {real, imag} */,
  {32'hc27d4eae, 32'hc231b2c2} /* (11, 29, 13) {real, imag} */,
  {32'hc125b563, 32'hc1aa4e6a} /* (11, 29, 12) {real, imag} */,
  {32'hc206a812, 32'h4195ad96} /* (11, 29, 11) {real, imag} */,
  {32'h42465da2, 32'hc1edbe04} /* (11, 29, 10) {real, imag} */,
  {32'hc1d7de8c, 32'h417b9dc4} /* (11, 29, 9) {real, imag} */,
  {32'hc1ffffce, 32'hc1dd7e6c} /* (11, 29, 8) {real, imag} */,
  {32'hc158b272, 32'hc27a85f4} /* (11, 29, 7) {real, imag} */,
  {32'h418a0b14, 32'h424bacec} /* (11, 29, 6) {real, imag} */,
  {32'hc3784552, 32'h41e64ce9} /* (11, 29, 5) {real, imag} */,
  {32'h43373972, 32'h429b6327} /* (11, 29, 4) {real, imag} */,
  {32'h4233475d, 32'hbfab3c50} /* (11, 29, 3) {real, imag} */,
  {32'hc4b8fc2c, 32'hc408e4b9} /* (11, 29, 2) {real, imag} */,
  {32'h459892e6, 32'h44b245c2} /* (11, 29, 1) {real, imag} */,
  {32'h45b01a21, 32'h00000000} /* (11, 29, 0) {real, imag} */,
  {32'h45a4369e, 32'hc4985aed} /* (11, 28, 31) {real, imag} */,
  {32'hc4d36833, 32'h43c6d004} /* (11, 28, 30) {real, imag} */,
  {32'h427e63ee, 32'h42f51838} /* (11, 28, 29) {real, imag} */,
  {32'h42afe1a6, 32'hc2ea9b94} /* (11, 28, 28) {real, imag} */,
  {32'hc3492f4c, 32'h429541fa} /* (11, 28, 27) {real, imag} */,
  {32'h40d17a5e, 32'h4255db24} /* (11, 28, 26) {real, imag} */,
  {32'h41a57227, 32'hc299eb31} /* (11, 28, 25) {real, imag} */,
  {32'hc31012c3, 32'h42362322} /* (11, 28, 24) {real, imag} */,
  {32'hc1f6e1dc, 32'h42df66c4} /* (11, 28, 23) {real, imag} */,
  {32'hc1c97f6e, 32'hc1a26a82} /* (11, 28, 22) {real, imag} */,
  {32'hc10ece18, 32'hc187efbd} /* (11, 28, 21) {real, imag} */,
  {32'h4296a614, 32'h4255c302} /* (11, 28, 20) {real, imag} */,
  {32'hc29b1e8e, 32'hc11cdf34} /* (11, 28, 19) {real, imag} */,
  {32'h41f0732e, 32'hc0e7a68c} /* (11, 28, 18) {real, imag} */,
  {32'h41ab9ca8, 32'hc2a7b7f0} /* (11, 28, 17) {real, imag} */,
  {32'hc218f0ca, 32'h00000000} /* (11, 28, 16) {real, imag} */,
  {32'h41ab9ca8, 32'h42a7b7f0} /* (11, 28, 15) {real, imag} */,
  {32'h41f0732e, 32'h40e7a68c} /* (11, 28, 14) {real, imag} */,
  {32'hc29b1e8e, 32'h411cdf34} /* (11, 28, 13) {real, imag} */,
  {32'h4296a614, 32'hc255c302} /* (11, 28, 12) {real, imag} */,
  {32'hc10ece18, 32'h4187efbd} /* (11, 28, 11) {real, imag} */,
  {32'hc1c97f6e, 32'h41a26a82} /* (11, 28, 10) {real, imag} */,
  {32'hc1f6e1dc, 32'hc2df66c4} /* (11, 28, 9) {real, imag} */,
  {32'hc31012c3, 32'hc2362322} /* (11, 28, 8) {real, imag} */,
  {32'h41a57227, 32'h4299eb31} /* (11, 28, 7) {real, imag} */,
  {32'h40d17a5e, 32'hc255db24} /* (11, 28, 6) {real, imag} */,
  {32'hc3492f4c, 32'hc29541fa} /* (11, 28, 5) {real, imag} */,
  {32'h42afe1a6, 32'h42ea9b94} /* (11, 28, 4) {real, imag} */,
  {32'h427e63ee, 32'hc2f51838} /* (11, 28, 3) {real, imag} */,
  {32'hc4d36833, 32'hc3c6d004} /* (11, 28, 2) {real, imag} */,
  {32'h45a4369e, 32'h44985aed} /* (11, 28, 1) {real, imag} */,
  {32'h45acf012, 32'h00000000} /* (11, 28, 0) {real, imag} */,
  {32'h45a8072f, 32'hc480ab34} /* (11, 27, 31) {real, imag} */,
  {32'hc4e9f8aa, 32'h4394683e} /* (11, 27, 30) {real, imag} */,
  {32'hc1d11656, 32'h42ef62ea} /* (11, 27, 29) {real, imag} */,
  {32'h431ed6a8, 32'hc3808ee0} /* (11, 27, 28) {real, imag} */,
  {32'hc317835e, 32'h419788bc} /* (11, 27, 27) {real, imag} */,
  {32'hc231ec7b, 32'h42928ee0} /* (11, 27, 26) {real, imag} */,
  {32'hc1008b68, 32'hc306941a} /* (11, 27, 25) {real, imag} */,
  {32'hc275da3e, 32'h424d9bc7} /* (11, 27, 24) {real, imag} */,
  {32'h408092d8, 32'h42c3ed70} /* (11, 27, 23) {real, imag} */,
  {32'h432d46a5, 32'h42837b2b} /* (11, 27, 22) {real, imag} */,
  {32'h4213e9ce, 32'hc0a09510} /* (11, 27, 21) {real, imag} */,
  {32'hc317fe92, 32'hc27e9b8e} /* (11, 27, 20) {real, imag} */,
  {32'hc271a93a, 32'h41ba16a8} /* (11, 27, 19) {real, imag} */,
  {32'hc267eaa2, 32'hc238b1cf} /* (11, 27, 18) {real, imag} */,
  {32'h423c8b57, 32'hc283584b} /* (11, 27, 17) {real, imag} */,
  {32'h4128104c, 32'h00000000} /* (11, 27, 16) {real, imag} */,
  {32'h423c8b57, 32'h4283584b} /* (11, 27, 15) {real, imag} */,
  {32'hc267eaa2, 32'h4238b1cf} /* (11, 27, 14) {real, imag} */,
  {32'hc271a93a, 32'hc1ba16a8} /* (11, 27, 13) {real, imag} */,
  {32'hc317fe92, 32'h427e9b8e} /* (11, 27, 12) {real, imag} */,
  {32'h4213e9ce, 32'h40a09510} /* (11, 27, 11) {real, imag} */,
  {32'h432d46a5, 32'hc2837b2b} /* (11, 27, 10) {real, imag} */,
  {32'h408092d8, 32'hc2c3ed70} /* (11, 27, 9) {real, imag} */,
  {32'hc275da3e, 32'hc24d9bc7} /* (11, 27, 8) {real, imag} */,
  {32'hc1008b68, 32'h4306941a} /* (11, 27, 7) {real, imag} */,
  {32'hc231ec7b, 32'hc2928ee0} /* (11, 27, 6) {real, imag} */,
  {32'hc317835e, 32'hc19788bc} /* (11, 27, 5) {real, imag} */,
  {32'h431ed6a8, 32'h43808ee0} /* (11, 27, 4) {real, imag} */,
  {32'hc1d11656, 32'hc2ef62ea} /* (11, 27, 3) {real, imag} */,
  {32'hc4e9f8aa, 32'hc394683e} /* (11, 27, 2) {real, imag} */,
  {32'h45a8072f, 32'h4480ab34} /* (11, 27, 1) {real, imag} */,
  {32'h45a9eb1e, 32'h00000000} /* (11, 27, 0) {real, imag} */,
  {32'h45a3bb95, 32'hc459615c} /* (11, 26, 31) {real, imag} */,
  {32'hc4e4ee89, 32'h43594b68} /* (11, 26, 30) {real, imag} */,
  {32'h421918da, 32'hc239dc5a} /* (11, 26, 29) {real, imag} */,
  {32'h4312cb89, 32'hc2ba22ac} /* (11, 26, 28) {real, imag} */,
  {32'hc30b3f12, 32'h40f53e80} /* (11, 26, 27) {real, imag} */,
  {32'hc2cbde0e, 32'h4284d911} /* (11, 26, 26) {real, imag} */,
  {32'h41e96ad0, 32'hc25f22ef} /* (11, 26, 25) {real, imag} */,
  {32'h418bc2cf, 32'h42890ba5} /* (11, 26, 24) {real, imag} */,
  {32'hbfe21570, 32'h42327a35} /* (11, 26, 23) {real, imag} */,
  {32'h410da4d4, 32'h42747bfe} /* (11, 26, 22) {real, imag} */,
  {32'h41c35e6c, 32'h42858859} /* (11, 26, 21) {real, imag} */,
  {32'h420a7c1a, 32'h41457661} /* (11, 26, 20) {real, imag} */,
  {32'h4299b736, 32'h419fdce0} /* (11, 26, 19) {real, imag} */,
  {32'h422d628e, 32'h40fe51f8} /* (11, 26, 18) {real, imag} */,
  {32'hbfc6fe00, 32'h40686520} /* (11, 26, 17) {real, imag} */,
  {32'h41054b01, 32'h00000000} /* (11, 26, 16) {real, imag} */,
  {32'hbfc6fe00, 32'hc0686520} /* (11, 26, 15) {real, imag} */,
  {32'h422d628e, 32'hc0fe51f8} /* (11, 26, 14) {real, imag} */,
  {32'h4299b736, 32'hc19fdce0} /* (11, 26, 13) {real, imag} */,
  {32'h420a7c1a, 32'hc1457661} /* (11, 26, 12) {real, imag} */,
  {32'h41c35e6c, 32'hc2858859} /* (11, 26, 11) {real, imag} */,
  {32'h410da4d4, 32'hc2747bfe} /* (11, 26, 10) {real, imag} */,
  {32'hbfe21570, 32'hc2327a35} /* (11, 26, 9) {real, imag} */,
  {32'h418bc2cf, 32'hc2890ba5} /* (11, 26, 8) {real, imag} */,
  {32'h41e96ad0, 32'h425f22ef} /* (11, 26, 7) {real, imag} */,
  {32'hc2cbde0e, 32'hc284d911} /* (11, 26, 6) {real, imag} */,
  {32'hc30b3f12, 32'hc0f53e80} /* (11, 26, 5) {real, imag} */,
  {32'h4312cb89, 32'h42ba22ac} /* (11, 26, 4) {real, imag} */,
  {32'h421918da, 32'h4239dc5a} /* (11, 26, 3) {real, imag} */,
  {32'hc4e4ee89, 32'hc3594b68} /* (11, 26, 2) {real, imag} */,
  {32'h45a3bb95, 32'h4459615c} /* (11, 26, 1) {real, imag} */,
  {32'h45a0d45a, 32'h00000000} /* (11, 26, 0) {real, imag} */,
  {32'h45992ebd, 32'hc40c8d9f} /* (11, 25, 31) {real, imag} */,
  {32'hc4e9af5e, 32'h436ffb28} /* (11, 25, 30) {real, imag} */,
  {32'hc2afa8e6, 32'h4289dbce} /* (11, 25, 29) {real, imag} */,
  {32'h42a6f63a, 32'hc3025fba} /* (11, 25, 28) {real, imag} */,
  {32'hc2f00b29, 32'h43615f36} /* (11, 25, 27) {real, imag} */,
  {32'hc36c8b17, 32'hc3207fbc} /* (11, 25, 26) {real, imag} */,
  {32'h42c97c9d, 32'h4250e0db} /* (11, 25, 25) {real, imag} */,
  {32'hc1933eaa, 32'h4284038f} /* (11, 25, 24) {real, imag} */,
  {32'h42d64bca, 32'h426b00aa} /* (11, 25, 23) {real, imag} */,
  {32'hc1d959ea, 32'hc272fff0} /* (11, 25, 22) {real, imag} */,
  {32'hc2af23d8, 32'hc1dbbca0} /* (11, 25, 21) {real, imag} */,
  {32'hc1c2a7ee, 32'h41382c03} /* (11, 25, 20) {real, imag} */,
  {32'h42658973, 32'h41d21afb} /* (11, 25, 19) {real, imag} */,
  {32'h42072c40, 32'hc27978e3} /* (11, 25, 18) {real, imag} */,
  {32'h41f9c750, 32'h41ec00a7} /* (11, 25, 17) {real, imag} */,
  {32'hc24897d8, 32'h00000000} /* (11, 25, 16) {real, imag} */,
  {32'h41f9c750, 32'hc1ec00a7} /* (11, 25, 15) {real, imag} */,
  {32'h42072c40, 32'h427978e3} /* (11, 25, 14) {real, imag} */,
  {32'h42658973, 32'hc1d21afb} /* (11, 25, 13) {real, imag} */,
  {32'hc1c2a7ee, 32'hc1382c03} /* (11, 25, 12) {real, imag} */,
  {32'hc2af23d8, 32'h41dbbca0} /* (11, 25, 11) {real, imag} */,
  {32'hc1d959ea, 32'h4272fff0} /* (11, 25, 10) {real, imag} */,
  {32'h42d64bca, 32'hc26b00aa} /* (11, 25, 9) {real, imag} */,
  {32'hc1933eaa, 32'hc284038f} /* (11, 25, 8) {real, imag} */,
  {32'h42c97c9d, 32'hc250e0db} /* (11, 25, 7) {real, imag} */,
  {32'hc36c8b17, 32'h43207fbc} /* (11, 25, 6) {real, imag} */,
  {32'hc2f00b29, 32'hc3615f36} /* (11, 25, 5) {real, imag} */,
  {32'h42a6f63a, 32'h43025fba} /* (11, 25, 4) {real, imag} */,
  {32'hc2afa8e6, 32'hc289dbce} /* (11, 25, 3) {real, imag} */,
  {32'hc4e9af5e, 32'hc36ffb28} /* (11, 25, 2) {real, imag} */,
  {32'h45992ebd, 32'h440c8d9f} /* (11, 25, 1) {real, imag} */,
  {32'h45921d2f, 32'h00000000} /* (11, 25, 0) {real, imag} */,
  {32'h45886e20, 32'hc33b7598} /* (11, 24, 31) {real, imag} */,
  {32'hc4d9014c, 32'h42a605b4} /* (11, 24, 30) {real, imag} */,
  {32'hc3196de2, 32'h42eee5f2} /* (11, 24, 29) {real, imag} */,
  {32'h432abec4, 32'hc2ec349c} /* (11, 24, 28) {real, imag} */,
  {32'hc385be13, 32'h435733ca} /* (11, 24, 27) {real, imag} */,
  {32'hc2dfb9e2, 32'hc2bb6a0a} /* (11, 24, 26) {real, imag} */,
  {32'h412b0804, 32'h42183ff6} /* (11, 24, 25) {real, imag} */,
  {32'hc28c2594, 32'hc2a710c4} /* (11, 24, 24) {real, imag} */,
  {32'h41b5ee20, 32'hc260b637} /* (11, 24, 23) {real, imag} */,
  {32'h412f4644, 32'hc2a5d554} /* (11, 24, 22) {real, imag} */,
  {32'hc2ba27a4, 32'h426d4d72} /* (11, 24, 21) {real, imag} */,
  {32'h4293b79e, 32'h42da0844} /* (11, 24, 20) {real, imag} */,
  {32'hc2737652, 32'hc1b53674} /* (11, 24, 19) {real, imag} */,
  {32'h42b087b6, 32'hc113bba8} /* (11, 24, 18) {real, imag} */,
  {32'hc252ee2a, 32'h41e003d2} /* (11, 24, 17) {real, imag} */,
  {32'hc22371bc, 32'h00000000} /* (11, 24, 16) {real, imag} */,
  {32'hc252ee2a, 32'hc1e003d2} /* (11, 24, 15) {real, imag} */,
  {32'h42b087b6, 32'h4113bba8} /* (11, 24, 14) {real, imag} */,
  {32'hc2737652, 32'h41b53674} /* (11, 24, 13) {real, imag} */,
  {32'h4293b79e, 32'hc2da0844} /* (11, 24, 12) {real, imag} */,
  {32'hc2ba27a4, 32'hc26d4d72} /* (11, 24, 11) {real, imag} */,
  {32'h412f4644, 32'h42a5d554} /* (11, 24, 10) {real, imag} */,
  {32'h41b5ee20, 32'h4260b637} /* (11, 24, 9) {real, imag} */,
  {32'hc28c2594, 32'h42a710c4} /* (11, 24, 8) {real, imag} */,
  {32'h412b0804, 32'hc2183ff6} /* (11, 24, 7) {real, imag} */,
  {32'hc2dfb9e2, 32'h42bb6a0a} /* (11, 24, 6) {real, imag} */,
  {32'hc385be13, 32'hc35733ca} /* (11, 24, 5) {real, imag} */,
  {32'h432abec4, 32'h42ec349c} /* (11, 24, 4) {real, imag} */,
  {32'hc3196de2, 32'hc2eee5f2} /* (11, 24, 3) {real, imag} */,
  {32'hc4d9014c, 32'hc2a605b4} /* (11, 24, 2) {real, imag} */,
  {32'h45886e20, 32'h433b7598} /* (11, 24, 1) {real, imag} */,
  {32'h457c5762, 32'h00000000} /* (11, 24, 0) {real, imag} */,
  {32'h4560f4ae, 32'hc2fc9778} /* (11, 23, 31) {real, imag} */,
  {32'hc4a1f1e1, 32'h426691e4} /* (11, 23, 30) {real, imag} */,
  {32'hc2b58568, 32'h428dcccd} /* (11, 23, 29) {real, imag} */,
  {32'h434bd4b8, 32'hc3086ec6} /* (11, 23, 28) {real, imag} */,
  {32'hc358ecee, 32'h432c3746} /* (11, 23, 27) {real, imag} */,
  {32'hc162a1e4, 32'hc2519c4b} /* (11, 23, 26) {real, imag} */,
  {32'h41f0f60c, 32'hc25d5cad} /* (11, 23, 25) {real, imag} */,
  {32'hc20a3671, 32'h422e763a} /* (11, 23, 24) {real, imag} */,
  {32'hc18ee8f2, 32'hc0bda1be} /* (11, 23, 23) {real, imag} */,
  {32'hc07eb010, 32'hc0e89370} /* (11, 23, 22) {real, imag} */,
  {32'h421d70ac, 32'h42f117da} /* (11, 23, 21) {real, imag} */,
  {32'hbea10500, 32'h41008c00} /* (11, 23, 20) {real, imag} */,
  {32'hc2842f6a, 32'h40309a20} /* (11, 23, 19) {real, imag} */,
  {32'h41b85313, 32'h41ed3d1e} /* (11, 23, 18) {real, imag} */,
  {32'hc1487a93, 32'h421254b2} /* (11, 23, 17) {real, imag} */,
  {32'hc20e7ff8, 32'h00000000} /* (11, 23, 16) {real, imag} */,
  {32'hc1487a93, 32'hc21254b2} /* (11, 23, 15) {real, imag} */,
  {32'h41b85313, 32'hc1ed3d1e} /* (11, 23, 14) {real, imag} */,
  {32'hc2842f6a, 32'hc0309a20} /* (11, 23, 13) {real, imag} */,
  {32'hbea10500, 32'hc1008c00} /* (11, 23, 12) {real, imag} */,
  {32'h421d70ac, 32'hc2f117da} /* (11, 23, 11) {real, imag} */,
  {32'hc07eb010, 32'h40e89370} /* (11, 23, 10) {real, imag} */,
  {32'hc18ee8f2, 32'h40bda1be} /* (11, 23, 9) {real, imag} */,
  {32'hc20a3671, 32'hc22e763a} /* (11, 23, 8) {real, imag} */,
  {32'h41f0f60c, 32'h425d5cad} /* (11, 23, 7) {real, imag} */,
  {32'hc162a1e4, 32'h42519c4b} /* (11, 23, 6) {real, imag} */,
  {32'hc358ecee, 32'hc32c3746} /* (11, 23, 5) {real, imag} */,
  {32'h434bd4b8, 32'h43086ec6} /* (11, 23, 4) {real, imag} */,
  {32'hc2b58568, 32'hc28dcccd} /* (11, 23, 3) {real, imag} */,
  {32'hc4a1f1e1, 32'hc26691e4} /* (11, 23, 2) {real, imag} */,
  {32'h4560f4ae, 32'h42fc9778} /* (11, 23, 1) {real, imag} */,
  {32'h4545cda9, 32'h00000000} /* (11, 23, 0) {real, imag} */,
  {32'h4519e123, 32'hc3359606} /* (11, 22, 31) {real, imag} */,
  {32'hc452d5e6, 32'h423bb2f4} /* (11, 22, 30) {real, imag} */,
  {32'hc00295b8, 32'h4154a4ee} /* (11, 22, 29) {real, imag} */,
  {32'h4398e5f4, 32'hc32131b9} /* (11, 22, 28) {real, imag} */,
  {32'hc347fbba, 32'h435c6774} /* (11, 22, 27) {real, imag} */,
  {32'hc267d6ef, 32'h42bdd8f0} /* (11, 22, 26) {real, imag} */,
  {32'h42d31df9, 32'hc1ff5538} /* (11, 22, 25) {real, imag} */,
  {32'hc2bf5ac4, 32'h431f56c7} /* (11, 22, 24) {real, imag} */,
  {32'h416c8953, 32'h41fed07c} /* (11, 22, 23) {real, imag} */,
  {32'hc1920760, 32'h4239cbe2} /* (11, 22, 22) {real, imag} */,
  {32'h42961812, 32'h42acb5a3} /* (11, 22, 21) {real, imag} */,
  {32'hc25ae8f6, 32'h41352ae4} /* (11, 22, 20) {real, imag} */,
  {32'h41b1c95a, 32'h42503266} /* (11, 22, 19) {real, imag} */,
  {32'hc22a0da0, 32'h41cc554b} /* (11, 22, 18) {real, imag} */,
  {32'h42037e89, 32'hc22c4c2b} /* (11, 22, 17) {real, imag} */,
  {32'h41de6b42, 32'h00000000} /* (11, 22, 16) {real, imag} */,
  {32'h42037e89, 32'h422c4c2b} /* (11, 22, 15) {real, imag} */,
  {32'hc22a0da0, 32'hc1cc554b} /* (11, 22, 14) {real, imag} */,
  {32'h41b1c95a, 32'hc2503266} /* (11, 22, 13) {real, imag} */,
  {32'hc25ae8f6, 32'hc1352ae4} /* (11, 22, 12) {real, imag} */,
  {32'h42961812, 32'hc2acb5a3} /* (11, 22, 11) {real, imag} */,
  {32'hc1920760, 32'hc239cbe2} /* (11, 22, 10) {real, imag} */,
  {32'h416c8953, 32'hc1fed07c} /* (11, 22, 9) {real, imag} */,
  {32'hc2bf5ac4, 32'hc31f56c7} /* (11, 22, 8) {real, imag} */,
  {32'h42d31df9, 32'h41ff5538} /* (11, 22, 7) {real, imag} */,
  {32'hc267d6ef, 32'hc2bdd8f0} /* (11, 22, 6) {real, imag} */,
  {32'hc347fbba, 32'hc35c6774} /* (11, 22, 5) {real, imag} */,
  {32'h4398e5f4, 32'h432131b9} /* (11, 22, 4) {real, imag} */,
  {32'hc00295b8, 32'hc154a4ee} /* (11, 22, 3) {real, imag} */,
  {32'hc452d5e6, 32'hc23bb2f4} /* (11, 22, 2) {real, imag} */,
  {32'h4519e123, 32'h43359606} /* (11, 22, 1) {real, imag} */,
  {32'h45019cb3, 32'h00000000} /* (11, 22, 0) {real, imag} */,
  {32'h445b784e, 32'hc2750a60} /* (11, 21, 31) {real, imag} */,
  {32'hc321b0e4, 32'hc28d0462} /* (11, 21, 30) {real, imag} */,
  {32'hc2d02d80, 32'h424092de} /* (11, 21, 29) {real, imag} */,
  {32'hc1b90fe6, 32'hc1c93eac} /* (11, 21, 28) {real, imag} */,
  {32'hc2f27622, 32'h428debb9} /* (11, 21, 27) {real, imag} */,
  {32'h422f0588, 32'h41ed9024} /* (11, 21, 26) {real, imag} */,
  {32'hc23292e0, 32'h43006249} /* (11, 21, 25) {real, imag} */,
  {32'h42b39ebb, 32'h428b8f8e} /* (11, 21, 24) {real, imag} */,
  {32'h4268daaa, 32'hc1d7d8d6} /* (11, 21, 23) {real, imag} */,
  {32'hc23c2add, 32'hc2ab4bf4} /* (11, 21, 22) {real, imag} */,
  {32'h3f269680, 32'h42635284} /* (11, 21, 21) {real, imag} */,
  {32'hc231d8e2, 32'h424ffa2b} /* (11, 21, 20) {real, imag} */,
  {32'hc21ed1fd, 32'hc15513fb} /* (11, 21, 19) {real, imag} */,
  {32'hc2934198, 32'h4282a30e} /* (11, 21, 18) {real, imag} */,
  {32'hc0f6d1c6, 32'hc00e03a8} /* (11, 21, 17) {real, imag} */,
  {32'hc15f0d54, 32'h00000000} /* (11, 21, 16) {real, imag} */,
  {32'hc0f6d1c6, 32'h400e03a8} /* (11, 21, 15) {real, imag} */,
  {32'hc2934198, 32'hc282a30e} /* (11, 21, 14) {real, imag} */,
  {32'hc21ed1fd, 32'h415513fb} /* (11, 21, 13) {real, imag} */,
  {32'hc231d8e2, 32'hc24ffa2b} /* (11, 21, 12) {real, imag} */,
  {32'h3f269680, 32'hc2635284} /* (11, 21, 11) {real, imag} */,
  {32'hc23c2add, 32'h42ab4bf4} /* (11, 21, 10) {real, imag} */,
  {32'h4268daaa, 32'h41d7d8d6} /* (11, 21, 9) {real, imag} */,
  {32'h42b39ebb, 32'hc28b8f8e} /* (11, 21, 8) {real, imag} */,
  {32'hc23292e0, 32'hc3006249} /* (11, 21, 7) {real, imag} */,
  {32'h422f0588, 32'hc1ed9024} /* (11, 21, 6) {real, imag} */,
  {32'hc2f27622, 32'hc28debb9} /* (11, 21, 5) {real, imag} */,
  {32'hc1b90fe6, 32'h41c93eac} /* (11, 21, 4) {real, imag} */,
  {32'hc2d02d80, 32'hc24092de} /* (11, 21, 3) {real, imag} */,
  {32'hc321b0e4, 32'h428d0462} /* (11, 21, 2) {real, imag} */,
  {32'h445b784e, 32'h42750a60} /* (11, 21, 1) {real, imag} */,
  {32'h44515a39, 32'h00000000} /* (11, 21, 0) {real, imag} */,
  {32'hc497f486, 32'h42f16e30} /* (11, 20, 31) {real, imag} */,
  {32'h441ce1a6, 32'hc3806376} /* (11, 20, 30) {real, imag} */,
  {32'hc33c2661, 32'h42225d5e} /* (11, 20, 29) {real, imag} */,
  {32'hc26a418c, 32'h42ce53a8} /* (11, 20, 28) {real, imag} */,
  {32'h42939b2b, 32'hc1605b9a} /* (11, 20, 27) {real, imag} */,
  {32'h42819af3, 32'h41f3ef22} /* (11, 20, 26) {real, imag} */,
  {32'hc19aace8, 32'hc2e6e443} /* (11, 20, 25) {real, imag} */,
  {32'h42dc91b0, 32'hc33552dc} /* (11, 20, 24) {real, imag} */,
  {32'h41be155b, 32'h421cb7df} /* (11, 20, 23) {real, imag} */,
  {32'h426a132b, 32'hc220c164} /* (11, 20, 22) {real, imag} */,
  {32'h42eae760, 32'hc1cd4016} /* (11, 20, 21) {real, imag} */,
  {32'hc1181001, 32'hc1f282ad} /* (11, 20, 20) {real, imag} */,
  {32'hc2b653d9, 32'h409283a4} /* (11, 20, 19) {real, imag} */,
  {32'h42436582, 32'hc12b6ba1} /* (11, 20, 18) {real, imag} */,
  {32'h40c31c60, 32'h3f353e60} /* (11, 20, 17) {real, imag} */,
  {32'hc146ff1c, 32'h00000000} /* (11, 20, 16) {real, imag} */,
  {32'h40c31c60, 32'hbf353e60} /* (11, 20, 15) {real, imag} */,
  {32'h42436582, 32'h412b6ba1} /* (11, 20, 14) {real, imag} */,
  {32'hc2b653d9, 32'hc09283a4} /* (11, 20, 13) {real, imag} */,
  {32'hc1181001, 32'h41f282ad} /* (11, 20, 12) {real, imag} */,
  {32'h42eae760, 32'h41cd4016} /* (11, 20, 11) {real, imag} */,
  {32'h426a132b, 32'h4220c164} /* (11, 20, 10) {real, imag} */,
  {32'h41be155b, 32'hc21cb7df} /* (11, 20, 9) {real, imag} */,
  {32'h42dc91b0, 32'h433552dc} /* (11, 20, 8) {real, imag} */,
  {32'hc19aace8, 32'h42e6e443} /* (11, 20, 7) {real, imag} */,
  {32'h42819af3, 32'hc1f3ef22} /* (11, 20, 6) {real, imag} */,
  {32'h42939b2b, 32'h41605b9a} /* (11, 20, 5) {real, imag} */,
  {32'hc26a418c, 32'hc2ce53a8} /* (11, 20, 4) {real, imag} */,
  {32'hc33c2661, 32'hc2225d5e} /* (11, 20, 3) {real, imag} */,
  {32'h441ce1a6, 32'h43806376} /* (11, 20, 2) {real, imag} */,
  {32'hc497f486, 32'hc2f16e30} /* (11, 20, 1) {real, imag} */,
  {32'hc42306cc, 32'h00000000} /* (11, 20, 0) {real, imag} */,
  {32'hc523dafd, 32'h439e8b70} /* (11, 19, 31) {real, imag} */,
  {32'h448ae62f, 32'hc3791277} /* (11, 19, 30) {real, imag} */,
  {32'hc2be5a37, 32'h4254ec4b} /* (11, 19, 29) {real, imag} */,
  {32'hc10f39a8, 32'hc1bf4b44} /* (11, 19, 28) {real, imag} */,
  {32'h431efa18, 32'h42b78bac} /* (11, 19, 27) {real, imag} */,
  {32'h42ed55c8, 32'h4206ae5e} /* (11, 19, 26) {real, imag} */,
  {32'hc187b0e9, 32'h41e8b5a1} /* (11, 19, 25) {real, imag} */,
  {32'h42d6c262, 32'hc32329c0} /* (11, 19, 24) {real, imag} */,
  {32'hc2c216a0, 32'h41857b8a} /* (11, 19, 23) {real, imag} */,
  {32'hc25dcc3a, 32'hc1c6c538} /* (11, 19, 22) {real, imag} */,
  {32'h4219aa6e, 32'hc29ab084} /* (11, 19, 21) {real, imag} */,
  {32'hc2d52d88, 32'hc2025308} /* (11, 19, 20) {real, imag} */,
  {32'h42100922, 32'h42e34a3e} /* (11, 19, 19) {real, imag} */,
  {32'hc173f230, 32'hc25847d5} /* (11, 19, 18) {real, imag} */,
  {32'h40baf51b, 32'hc10e333c} /* (11, 19, 17) {real, imag} */,
  {32'hc27f22a4, 32'h00000000} /* (11, 19, 16) {real, imag} */,
  {32'h40baf51b, 32'h410e333c} /* (11, 19, 15) {real, imag} */,
  {32'hc173f230, 32'h425847d5} /* (11, 19, 14) {real, imag} */,
  {32'h42100922, 32'hc2e34a3e} /* (11, 19, 13) {real, imag} */,
  {32'hc2d52d88, 32'h42025308} /* (11, 19, 12) {real, imag} */,
  {32'h4219aa6e, 32'h429ab084} /* (11, 19, 11) {real, imag} */,
  {32'hc25dcc3a, 32'h41c6c538} /* (11, 19, 10) {real, imag} */,
  {32'hc2c216a0, 32'hc1857b8a} /* (11, 19, 9) {real, imag} */,
  {32'h42d6c262, 32'h432329c0} /* (11, 19, 8) {real, imag} */,
  {32'hc187b0e9, 32'hc1e8b5a1} /* (11, 19, 7) {real, imag} */,
  {32'h42ed55c8, 32'hc206ae5e} /* (11, 19, 6) {real, imag} */,
  {32'h431efa18, 32'hc2b78bac} /* (11, 19, 5) {real, imag} */,
  {32'hc10f39a8, 32'h41bf4b44} /* (11, 19, 4) {real, imag} */,
  {32'hc2be5a37, 32'hc254ec4b} /* (11, 19, 3) {real, imag} */,
  {32'h448ae62f, 32'h43791277} /* (11, 19, 2) {real, imag} */,
  {32'hc523dafd, 32'hc39e8b70} /* (11, 19, 1) {real, imag} */,
  {32'hc4e2e5e6, 32'h00000000} /* (11, 19, 0) {real, imag} */,
  {32'hc558d576, 32'h43d063c0} /* (11, 18, 31) {real, imag} */,
  {32'h44a8962e, 32'hc35292f3} /* (11, 18, 30) {real, imag} */,
  {32'h428582f5, 32'h42a98f3b} /* (11, 18, 29) {real, imag} */,
  {32'hc2c3e468, 32'h4318c550} /* (11, 18, 28) {real, imag} */,
  {32'h4340b5c6, 32'h40fcd790} /* (11, 18, 27) {real, imag} */,
  {32'hc19b3285, 32'hc30407cf} /* (11, 18, 26) {real, imag} */,
  {32'h42224324, 32'h41813c08} /* (11, 18, 25) {real, imag} */,
  {32'h43199f30, 32'hc1e41bdc} /* (11, 18, 24) {real, imag} */,
  {32'hc2628eda, 32'h4069c338} /* (11, 18, 23) {real, imag} */,
  {32'h41d4c5b2, 32'hc2621f2e} /* (11, 18, 22) {real, imag} */,
  {32'h4286874e, 32'h4212f798} /* (11, 18, 21) {real, imag} */,
  {32'h42957c14, 32'h41c2d669} /* (11, 18, 20) {real, imag} */,
  {32'h408891c8, 32'h420f95a3} /* (11, 18, 19) {real, imag} */,
  {32'hc2c0189f, 32'hc1c22a18} /* (11, 18, 18) {real, imag} */,
  {32'h42843177, 32'hc19f242d} /* (11, 18, 17) {real, imag} */,
  {32'hc2819754, 32'h00000000} /* (11, 18, 16) {real, imag} */,
  {32'h42843177, 32'h419f242d} /* (11, 18, 15) {real, imag} */,
  {32'hc2c0189f, 32'h41c22a18} /* (11, 18, 14) {real, imag} */,
  {32'h408891c8, 32'hc20f95a3} /* (11, 18, 13) {real, imag} */,
  {32'h42957c14, 32'hc1c2d669} /* (11, 18, 12) {real, imag} */,
  {32'h4286874e, 32'hc212f798} /* (11, 18, 11) {real, imag} */,
  {32'h41d4c5b2, 32'h42621f2e} /* (11, 18, 10) {real, imag} */,
  {32'hc2628eda, 32'hc069c338} /* (11, 18, 9) {real, imag} */,
  {32'h43199f30, 32'h41e41bdc} /* (11, 18, 8) {real, imag} */,
  {32'h42224324, 32'hc1813c08} /* (11, 18, 7) {real, imag} */,
  {32'hc19b3285, 32'h430407cf} /* (11, 18, 6) {real, imag} */,
  {32'h4340b5c6, 32'hc0fcd790} /* (11, 18, 5) {real, imag} */,
  {32'hc2c3e468, 32'hc318c550} /* (11, 18, 4) {real, imag} */,
  {32'h428582f5, 32'hc2a98f3b} /* (11, 18, 3) {real, imag} */,
  {32'h44a8962e, 32'h435292f3} /* (11, 18, 2) {real, imag} */,
  {32'hc558d576, 32'hc3d063c0} /* (11, 18, 1) {real, imag} */,
  {32'hc52e3a92, 32'h00000000} /* (11, 18, 0) {real, imag} */,
  {32'hc58204aa, 32'h43ae0266} /* (11, 17, 31) {real, imag} */,
  {32'h44c712cf, 32'hc3dfce92} /* (11, 17, 30) {real, imag} */,
  {32'h42e0e99f, 32'hc30d9df8} /* (11, 17, 29) {real, imag} */,
  {32'hc26177b8, 32'h42be2b0d} /* (11, 17, 28) {real, imag} */,
  {32'h43b05931, 32'hc2a88e10} /* (11, 17, 27) {real, imag} */,
  {32'hc2910758, 32'hc2b3dc54} /* (11, 17, 26) {real, imag} */,
  {32'h42c7d0b4, 32'h3fc0f700} /* (11, 17, 25) {real, imag} */,
  {32'h421b2752, 32'h427de0e1} /* (11, 17, 24) {real, imag} */,
  {32'h418012fc, 32'h42cbe230} /* (11, 17, 23) {real, imag} */,
  {32'hc2ec5230, 32'hc1dc4962} /* (11, 17, 22) {real, imag} */,
  {32'hc2569445, 32'hc1284dbb} /* (11, 17, 21) {real, imag} */,
  {32'h3f389120, 32'hc0c31a4c} /* (11, 17, 20) {real, imag} */,
  {32'h41f40b75, 32'hc27c3ef5} /* (11, 17, 19) {real, imag} */,
  {32'h4194e3e4, 32'hc202040a} /* (11, 17, 18) {real, imag} */,
  {32'hc239a7f8, 32'h4288922d} /* (11, 17, 17) {real, imag} */,
  {32'h4220c96f, 32'h00000000} /* (11, 17, 16) {real, imag} */,
  {32'hc239a7f8, 32'hc288922d} /* (11, 17, 15) {real, imag} */,
  {32'h4194e3e4, 32'h4202040a} /* (11, 17, 14) {real, imag} */,
  {32'h41f40b75, 32'h427c3ef5} /* (11, 17, 13) {real, imag} */,
  {32'h3f389120, 32'h40c31a4c} /* (11, 17, 12) {real, imag} */,
  {32'hc2569445, 32'h41284dbb} /* (11, 17, 11) {real, imag} */,
  {32'hc2ec5230, 32'h41dc4962} /* (11, 17, 10) {real, imag} */,
  {32'h418012fc, 32'hc2cbe230} /* (11, 17, 9) {real, imag} */,
  {32'h421b2752, 32'hc27de0e1} /* (11, 17, 8) {real, imag} */,
  {32'h42c7d0b4, 32'hbfc0f700} /* (11, 17, 7) {real, imag} */,
  {32'hc2910758, 32'h42b3dc54} /* (11, 17, 6) {real, imag} */,
  {32'h43b05931, 32'h42a88e10} /* (11, 17, 5) {real, imag} */,
  {32'hc26177b8, 32'hc2be2b0d} /* (11, 17, 4) {real, imag} */,
  {32'h42e0e99f, 32'h430d9df8} /* (11, 17, 3) {real, imag} */,
  {32'h44c712cf, 32'h43dfce92} /* (11, 17, 2) {real, imag} */,
  {32'hc58204aa, 32'hc3ae0266} /* (11, 17, 1) {real, imag} */,
  {32'hc5471511, 32'h00000000} /* (11, 17, 0) {real, imag} */,
  {32'hc58bcc0c, 32'h43ab2150} /* (11, 16, 31) {real, imag} */,
  {32'h44cdffc1, 32'hc399da60} /* (11, 16, 30) {real, imag} */,
  {32'h419eb15c, 32'h407b0360} /* (11, 16, 29) {real, imag} */,
  {32'hc32bb718, 32'hc2965800} /* (11, 16, 28) {real, imag} */,
  {32'h43a01792, 32'hc30f6c24} /* (11, 16, 27) {real, imag} */,
  {32'h429df442, 32'h4224a6e0} /* (11, 16, 26) {real, imag} */,
  {32'hc0a61d78, 32'h422e0100} /* (11, 16, 25) {real, imag} */,
  {32'h409b4eac, 32'h421e2b0a} /* (11, 16, 24) {real, imag} */,
  {32'hc1cd9e07, 32'h42c1cc32} /* (11, 16, 23) {real, imag} */,
  {32'h429a08bf, 32'h41ae4f03} /* (11, 16, 22) {real, imag} */,
  {32'hc0ff64d8, 32'hc246e4d8} /* (11, 16, 21) {real, imag} */,
  {32'hc1740d08, 32'h422723a6} /* (11, 16, 20) {real, imag} */,
  {32'hc207d0ee, 32'hc2618b5c} /* (11, 16, 19) {real, imag} */,
  {32'hc09fb48e, 32'hc2f58fc6} /* (11, 16, 18) {real, imag} */,
  {32'hc02afae8, 32'hc1cc7937} /* (11, 16, 17) {real, imag} */,
  {32'h42159ddd, 32'h00000000} /* (11, 16, 16) {real, imag} */,
  {32'hc02afae8, 32'h41cc7937} /* (11, 16, 15) {real, imag} */,
  {32'hc09fb48e, 32'h42f58fc6} /* (11, 16, 14) {real, imag} */,
  {32'hc207d0ee, 32'h42618b5c} /* (11, 16, 13) {real, imag} */,
  {32'hc1740d08, 32'hc22723a6} /* (11, 16, 12) {real, imag} */,
  {32'hc0ff64d8, 32'h4246e4d8} /* (11, 16, 11) {real, imag} */,
  {32'h429a08bf, 32'hc1ae4f03} /* (11, 16, 10) {real, imag} */,
  {32'hc1cd9e07, 32'hc2c1cc32} /* (11, 16, 9) {real, imag} */,
  {32'h409b4eac, 32'hc21e2b0a} /* (11, 16, 8) {real, imag} */,
  {32'hc0a61d78, 32'hc22e0100} /* (11, 16, 7) {real, imag} */,
  {32'h429df442, 32'hc224a6e0} /* (11, 16, 6) {real, imag} */,
  {32'h43a01792, 32'h430f6c24} /* (11, 16, 5) {real, imag} */,
  {32'hc32bb718, 32'h42965800} /* (11, 16, 4) {real, imag} */,
  {32'h419eb15c, 32'hc07b0360} /* (11, 16, 3) {real, imag} */,
  {32'h44cdffc1, 32'h4399da60} /* (11, 16, 2) {real, imag} */,
  {32'hc58bcc0c, 32'hc3ab2150} /* (11, 16, 1) {real, imag} */,
  {32'hc558eb8f, 32'h00000000} /* (11, 16, 0) {real, imag} */,
  {32'hc58cce12, 32'h4362aa54} /* (11, 15, 31) {real, imag} */,
  {32'h44c6299f, 32'hc32c3f94} /* (11, 15, 30) {real, imag} */,
  {32'h42c5ac13, 32'h4292cc54} /* (11, 15, 29) {real, imag} */,
  {32'hc3752226, 32'hc211542e} /* (11, 15, 28) {real, imag} */,
  {32'h4317c066, 32'hc20d39c0} /* (11, 15, 27) {real, imag} */,
  {32'h433add4e, 32'hc22eb4dc} /* (11, 15, 26) {real, imag} */,
  {32'hc2a54b72, 32'h4099c940} /* (11, 15, 25) {real, imag} */,
  {32'h4270b9a6, 32'hc03eb9f0} /* (11, 15, 24) {real, imag} */,
  {32'h42512e5c, 32'hc2513c71} /* (11, 15, 23) {real, imag} */,
  {32'hc2b2b3fa, 32'hc2b91586} /* (11, 15, 22) {real, imag} */,
  {32'hc0a13068, 32'hc109d823} /* (11, 15, 21) {real, imag} */,
  {32'h4215dd8a, 32'hc2213774} /* (11, 15, 20) {real, imag} */,
  {32'hc24fae2a, 32'h4214daa3} /* (11, 15, 19) {real, imag} */,
  {32'hc2283d32, 32'hc1e03aa5} /* (11, 15, 18) {real, imag} */,
  {32'h414408a2, 32'hc1bfeddf} /* (11, 15, 17) {real, imag} */,
  {32'hc27aa283, 32'h00000000} /* (11, 15, 16) {real, imag} */,
  {32'h414408a2, 32'h41bfeddf} /* (11, 15, 15) {real, imag} */,
  {32'hc2283d32, 32'h41e03aa5} /* (11, 15, 14) {real, imag} */,
  {32'hc24fae2a, 32'hc214daa3} /* (11, 15, 13) {real, imag} */,
  {32'h4215dd8a, 32'h42213774} /* (11, 15, 12) {real, imag} */,
  {32'hc0a13068, 32'h4109d823} /* (11, 15, 11) {real, imag} */,
  {32'hc2b2b3fa, 32'h42b91586} /* (11, 15, 10) {real, imag} */,
  {32'h42512e5c, 32'h42513c71} /* (11, 15, 9) {real, imag} */,
  {32'h4270b9a6, 32'h403eb9f0} /* (11, 15, 8) {real, imag} */,
  {32'hc2a54b72, 32'hc099c940} /* (11, 15, 7) {real, imag} */,
  {32'h433add4e, 32'h422eb4dc} /* (11, 15, 6) {real, imag} */,
  {32'h4317c066, 32'h420d39c0} /* (11, 15, 5) {real, imag} */,
  {32'hc3752226, 32'h4211542e} /* (11, 15, 4) {real, imag} */,
  {32'h42c5ac13, 32'hc292cc54} /* (11, 15, 3) {real, imag} */,
  {32'h44c6299f, 32'h432c3f94} /* (11, 15, 2) {real, imag} */,
  {32'hc58cce12, 32'hc362aa54} /* (11, 15, 1) {real, imag} */,
  {32'hc559130b, 32'h00000000} /* (11, 15, 0) {real, imag} */,
  {32'hc586113b, 32'h43be95d0} /* (11, 14, 31) {real, imag} */,
  {32'h44b04dfa, 32'hc3953202} /* (11, 14, 30) {real, imag} */,
  {32'hc119e8d8, 32'h42d59d15} /* (11, 14, 29) {real, imag} */,
  {32'hc3879ff8, 32'h4305d612} /* (11, 14, 28) {real, imag} */,
  {32'h43780562, 32'hc3112d46} /* (11, 14, 27) {real, imag} */,
  {32'h420e1a22, 32'hc1b992f0} /* (11, 14, 26) {real, imag} */,
  {32'h42ad7235, 32'h423cf52c} /* (11, 14, 25) {real, imag} */,
  {32'h42b4adea, 32'hc2d13757} /* (11, 14, 24) {real, imag} */,
  {32'hc1c39b8c, 32'hc18a6fd7} /* (11, 14, 23) {real, imag} */,
  {32'hc2722825, 32'hc2f40817} /* (11, 14, 22) {real, imag} */,
  {32'h3facaae0, 32'hc2bf76ee} /* (11, 14, 21) {real, imag} */,
  {32'hc2eef614, 32'h41c38f9b} /* (11, 14, 20) {real, imag} */,
  {32'h42afa92e, 32'hc1400494} /* (11, 14, 19) {real, imag} */,
  {32'hc19c6054, 32'h3fbd82d8} /* (11, 14, 18) {real, imag} */,
  {32'hc2af5eff, 32'hc085accc} /* (11, 14, 17) {real, imag} */,
  {32'h4251758a, 32'h00000000} /* (11, 14, 16) {real, imag} */,
  {32'hc2af5eff, 32'h4085accc} /* (11, 14, 15) {real, imag} */,
  {32'hc19c6054, 32'hbfbd82d8} /* (11, 14, 14) {real, imag} */,
  {32'h42afa92e, 32'h41400494} /* (11, 14, 13) {real, imag} */,
  {32'hc2eef614, 32'hc1c38f9b} /* (11, 14, 12) {real, imag} */,
  {32'h3facaae0, 32'h42bf76ee} /* (11, 14, 11) {real, imag} */,
  {32'hc2722825, 32'h42f40817} /* (11, 14, 10) {real, imag} */,
  {32'hc1c39b8c, 32'h418a6fd7} /* (11, 14, 9) {real, imag} */,
  {32'h42b4adea, 32'h42d13757} /* (11, 14, 8) {real, imag} */,
  {32'h42ad7235, 32'hc23cf52c} /* (11, 14, 7) {real, imag} */,
  {32'h420e1a22, 32'h41b992f0} /* (11, 14, 6) {real, imag} */,
  {32'h43780562, 32'h43112d46} /* (11, 14, 5) {real, imag} */,
  {32'hc3879ff8, 32'hc305d612} /* (11, 14, 4) {real, imag} */,
  {32'hc119e8d8, 32'hc2d59d15} /* (11, 14, 3) {real, imag} */,
  {32'h44b04dfa, 32'h43953202} /* (11, 14, 2) {real, imag} */,
  {32'hc586113b, 32'hc3be95d0} /* (11, 14, 1) {real, imag} */,
  {32'hc5448036, 32'h00000000} /* (11, 14, 0) {real, imag} */,
  {32'hc5650067, 32'h438ebf40} /* (11, 13, 31) {real, imag} */,
  {32'h44a62355, 32'hc2ef1812} /* (11, 13, 30) {real, imag} */,
  {32'hc2cffc1d, 32'h42432759} /* (11, 13, 29) {real, imag} */,
  {32'hc33d9ae6, 32'h43829d53} /* (11, 13, 28) {real, imag} */,
  {32'h42d7b830, 32'hc263f1af} /* (11, 13, 27) {real, imag} */,
  {32'hc09b2cb0, 32'h4208bab0} /* (11, 13, 26) {real, imag} */,
  {32'h4234b468, 32'h41c568fb} /* (11, 13, 25) {real, imag} */,
  {32'h42f58d76, 32'hc2d365eb} /* (11, 13, 24) {real, imag} */,
  {32'h40e52318, 32'h42b76640} /* (11, 13, 23) {real, imag} */,
  {32'h40e02ae4, 32'h42514d54} /* (11, 13, 22) {real, imag} */,
  {32'h414c5058, 32'hc11a8e2c} /* (11, 13, 21) {real, imag} */,
  {32'h422e9f78, 32'hc2cd8f38} /* (11, 13, 20) {real, imag} */,
  {32'h4248fa28, 32'hc327c4f5} /* (11, 13, 19) {real, imag} */,
  {32'hc1f43954, 32'hc25e4397} /* (11, 13, 18) {real, imag} */,
  {32'hc1820dfe, 32'h425f04b3} /* (11, 13, 17) {real, imag} */,
  {32'hc2b12b56, 32'h00000000} /* (11, 13, 16) {real, imag} */,
  {32'hc1820dfe, 32'hc25f04b3} /* (11, 13, 15) {real, imag} */,
  {32'hc1f43954, 32'h425e4397} /* (11, 13, 14) {real, imag} */,
  {32'h4248fa28, 32'h4327c4f5} /* (11, 13, 13) {real, imag} */,
  {32'h422e9f78, 32'h42cd8f38} /* (11, 13, 12) {real, imag} */,
  {32'h414c5058, 32'h411a8e2c} /* (11, 13, 11) {real, imag} */,
  {32'h40e02ae4, 32'hc2514d54} /* (11, 13, 10) {real, imag} */,
  {32'h40e52318, 32'hc2b76640} /* (11, 13, 9) {real, imag} */,
  {32'h42f58d76, 32'h42d365eb} /* (11, 13, 8) {real, imag} */,
  {32'h4234b468, 32'hc1c568fb} /* (11, 13, 7) {real, imag} */,
  {32'hc09b2cb0, 32'hc208bab0} /* (11, 13, 6) {real, imag} */,
  {32'h42d7b830, 32'h4263f1af} /* (11, 13, 5) {real, imag} */,
  {32'hc33d9ae6, 32'hc3829d53} /* (11, 13, 4) {real, imag} */,
  {32'hc2cffc1d, 32'hc2432759} /* (11, 13, 3) {real, imag} */,
  {32'h44a62355, 32'h42ef1812} /* (11, 13, 2) {real, imag} */,
  {32'hc5650067, 32'hc38ebf40} /* (11, 13, 1) {real, imag} */,
  {32'hc51b06ad, 32'h00000000} /* (11, 13, 0) {real, imag} */,
  {32'hc528de1d, 32'hc272cbe0} /* (11, 12, 31) {real, imag} */,
  {32'h448e2ead, 32'hc31a29cc} /* (11, 12, 30) {real, imag} */,
  {32'hc33e367f, 32'hc1d2fc24} /* (11, 12, 29) {real, imag} */,
  {32'hc27412f4, 32'h43298bec} /* (11, 12, 28) {real, imag} */,
  {32'h431f79fc, 32'hc1a0ea65} /* (11, 12, 27) {real, imag} */,
  {32'hc221888e, 32'hc0c1d890} /* (11, 12, 26) {real, imag} */,
  {32'hc2059e29, 32'hc2a1627d} /* (11, 12, 25) {real, imag} */,
  {32'h41e027be, 32'hc1c37eb4} /* (11, 12, 24) {real, imag} */,
  {32'h41bb8a55, 32'h419b7c8a} /* (11, 12, 23) {real, imag} */,
  {32'h42023d5f, 32'hc1c813a9} /* (11, 12, 22) {real, imag} */,
  {32'h422480c0, 32'hc005b5cc} /* (11, 12, 21) {real, imag} */,
  {32'h401cff4c, 32'h41a0dab5} /* (11, 12, 20) {real, imag} */,
  {32'h4254e6fe, 32'hc1565a68} /* (11, 12, 19) {real, imag} */,
  {32'h425ff536, 32'hc0dd226e} /* (11, 12, 18) {real, imag} */,
  {32'hc21efff8, 32'h423ec45a} /* (11, 12, 17) {real, imag} */,
  {32'h42000db9, 32'h00000000} /* (11, 12, 16) {real, imag} */,
  {32'hc21efff8, 32'hc23ec45a} /* (11, 12, 15) {real, imag} */,
  {32'h425ff536, 32'h40dd226e} /* (11, 12, 14) {real, imag} */,
  {32'h4254e6fe, 32'h41565a68} /* (11, 12, 13) {real, imag} */,
  {32'h401cff4c, 32'hc1a0dab5} /* (11, 12, 12) {real, imag} */,
  {32'h422480c0, 32'h4005b5cc} /* (11, 12, 11) {real, imag} */,
  {32'h42023d5f, 32'h41c813a9} /* (11, 12, 10) {real, imag} */,
  {32'h41bb8a55, 32'hc19b7c8a} /* (11, 12, 9) {real, imag} */,
  {32'h41e027be, 32'h41c37eb4} /* (11, 12, 8) {real, imag} */,
  {32'hc2059e29, 32'h42a1627d} /* (11, 12, 7) {real, imag} */,
  {32'hc221888e, 32'h40c1d890} /* (11, 12, 6) {real, imag} */,
  {32'h431f79fc, 32'h41a0ea65} /* (11, 12, 5) {real, imag} */,
  {32'hc27412f4, 32'hc3298bec} /* (11, 12, 4) {real, imag} */,
  {32'hc33e367f, 32'h41d2fc24} /* (11, 12, 3) {real, imag} */,
  {32'h448e2ead, 32'h431a29cc} /* (11, 12, 2) {real, imag} */,
  {32'hc528de1d, 32'h4272cbe0} /* (11, 12, 1) {real, imag} */,
  {32'hc4bd667a, 32'h00000000} /* (11, 12, 0) {real, imag} */,
  {32'hc4bb034f, 32'hc376b2b8} /* (11, 11, 31) {real, imag} */,
  {32'h442dace9, 32'hc2f1bb16} /* (11, 11, 30) {real, imag} */,
  {32'hc2acd6ca, 32'hc27b9c92} /* (11, 11, 29) {real, imag} */,
  {32'hc2f5c60e, 32'h428c6571} /* (11, 11, 28) {real, imag} */,
  {32'h42c8ecd2, 32'h42238392} /* (11, 11, 27) {real, imag} */,
  {32'h4338356c, 32'h421c427c} /* (11, 11, 26) {real, imag} */,
  {32'h40471f78, 32'h417c4254} /* (11, 11, 25) {real, imag} */,
  {32'h4274a7de, 32'h428a6a5a} /* (11, 11, 24) {real, imag} */,
  {32'hc30ff10e, 32'h4288d07c} /* (11, 11, 23) {real, imag} */,
  {32'h42f43b52, 32'hc289fc02} /* (11, 11, 22) {real, imag} */,
  {32'hc232be95, 32'hc258e664} /* (11, 11, 21) {real, imag} */,
  {32'h4185da85, 32'hc1d9d3b2} /* (11, 11, 20) {real, imag} */,
  {32'hc1d6bebe, 32'hc1a7ac50} /* (11, 11, 19) {real, imag} */,
  {32'h42aba90c, 32'h421a7c1a} /* (11, 11, 18) {real, imag} */,
  {32'hc1abadf2, 32'hc1a5cc99} /* (11, 11, 17) {real, imag} */,
  {32'h4288e08a, 32'h00000000} /* (11, 11, 16) {real, imag} */,
  {32'hc1abadf2, 32'h41a5cc99} /* (11, 11, 15) {real, imag} */,
  {32'h42aba90c, 32'hc21a7c1a} /* (11, 11, 14) {real, imag} */,
  {32'hc1d6bebe, 32'h41a7ac50} /* (11, 11, 13) {real, imag} */,
  {32'h4185da85, 32'h41d9d3b2} /* (11, 11, 12) {real, imag} */,
  {32'hc232be95, 32'h4258e664} /* (11, 11, 11) {real, imag} */,
  {32'h42f43b52, 32'h4289fc02} /* (11, 11, 10) {real, imag} */,
  {32'hc30ff10e, 32'hc288d07c} /* (11, 11, 9) {real, imag} */,
  {32'h4274a7de, 32'hc28a6a5a} /* (11, 11, 8) {real, imag} */,
  {32'h40471f78, 32'hc17c4254} /* (11, 11, 7) {real, imag} */,
  {32'h4338356c, 32'hc21c427c} /* (11, 11, 6) {real, imag} */,
  {32'h42c8ecd2, 32'hc2238392} /* (11, 11, 5) {real, imag} */,
  {32'hc2f5c60e, 32'hc28c6571} /* (11, 11, 4) {real, imag} */,
  {32'hc2acd6ca, 32'h427b9c92} /* (11, 11, 3) {real, imag} */,
  {32'h442dace9, 32'h42f1bb16} /* (11, 11, 2) {real, imag} */,
  {32'hc4bb034f, 32'h4376b2b8} /* (11, 11, 1) {real, imag} */,
  {32'hc39dfa72, 32'h00000000} /* (11, 11, 0) {real, imag} */,
  {32'h43d6abf8, 32'hc42c8c28} /* (11, 10, 31) {real, imag} */,
  {32'hc3960b07, 32'h432e397d} /* (11, 10, 30) {real, imag} */,
  {32'h418bf029, 32'hc2802946} /* (11, 10, 29) {real, imag} */,
  {32'hc21beabc, 32'hc37e30d7} /* (11, 10, 28) {real, imag} */,
  {32'hc1dd0204, 32'h43281fb8} /* (11, 10, 27) {real, imag} */,
  {32'h431bee4f, 32'hc15e4ad4} /* (11, 10, 26) {real, imag} */,
  {32'hc1164078, 32'h41cdbc5c} /* (11, 10, 25) {real, imag} */,
  {32'h415b0d94, 32'h428a219e} /* (11, 10, 24) {real, imag} */,
  {32'h4210760a, 32'h413ddd5b} /* (11, 10, 23) {real, imag} */,
  {32'hc0ec0c10, 32'h40568700} /* (11, 10, 22) {real, imag} */,
  {32'hc283cb38, 32'h42da94f5} /* (11, 10, 21) {real, imag} */,
  {32'hc25852fa, 32'h42a1f98a} /* (11, 10, 20) {real, imag} */,
  {32'hc22f2f87, 32'hc1790da8} /* (11, 10, 19) {real, imag} */,
  {32'h42982a38, 32'hc1ca535b} /* (11, 10, 18) {real, imag} */,
  {32'hc137abb4, 32'h41a45dfe} /* (11, 10, 17) {real, imag} */,
  {32'hc2829e62, 32'h00000000} /* (11, 10, 16) {real, imag} */,
  {32'hc137abb4, 32'hc1a45dfe} /* (11, 10, 15) {real, imag} */,
  {32'h42982a38, 32'h41ca535b} /* (11, 10, 14) {real, imag} */,
  {32'hc22f2f87, 32'h41790da8} /* (11, 10, 13) {real, imag} */,
  {32'hc25852fa, 32'hc2a1f98a} /* (11, 10, 12) {real, imag} */,
  {32'hc283cb38, 32'hc2da94f5} /* (11, 10, 11) {real, imag} */,
  {32'hc0ec0c10, 32'hc0568700} /* (11, 10, 10) {real, imag} */,
  {32'h4210760a, 32'hc13ddd5b} /* (11, 10, 9) {real, imag} */,
  {32'h415b0d94, 32'hc28a219e} /* (11, 10, 8) {real, imag} */,
  {32'hc1164078, 32'hc1cdbc5c} /* (11, 10, 7) {real, imag} */,
  {32'h431bee4f, 32'h415e4ad4} /* (11, 10, 6) {real, imag} */,
  {32'hc1dd0204, 32'hc3281fb8} /* (11, 10, 5) {real, imag} */,
  {32'hc21beabc, 32'h437e30d7} /* (11, 10, 4) {real, imag} */,
  {32'h418bf029, 32'h42802946} /* (11, 10, 3) {real, imag} */,
  {32'hc3960b07, 32'hc32e397d} /* (11, 10, 2) {real, imag} */,
  {32'h43d6abf8, 32'h442c8c28} /* (11, 10, 1) {real, imag} */,
  {32'h44b08b26, 32'h00000000} /* (11, 10, 0) {real, imag} */,
  {32'h44e5fbec, 32'hc4856cca} /* (11, 9, 31) {real, imag} */,
  {32'hc44e1142, 32'h439a51d4} /* (11, 9, 30) {real, imag} */,
  {32'hc2a89b66, 32'hc334ee74} /* (11, 9, 29) {real, imag} */,
  {32'h41c023e4, 32'hc2d756eb} /* (11, 9, 28) {real, imag} */,
  {32'hc2cb68b0, 32'h432ee31e} /* (11, 9, 27) {real, imag} */,
  {32'hc27fedb1, 32'h42aa8596} /* (11, 9, 26) {real, imag} */,
  {32'h4227a76c, 32'hc1b9c792} /* (11, 9, 25) {real, imag} */,
  {32'hc24db223, 32'hbf3d5ba0} /* (11, 9, 24) {real, imag} */,
  {32'h42bcbf9e, 32'hc1c90fa4} /* (11, 9, 23) {real, imag} */,
  {32'h429e5754, 32'h42a54814} /* (11, 9, 22) {real, imag} */,
  {32'h4246375a, 32'h41d90570} /* (11, 9, 21) {real, imag} */,
  {32'hc2779c3c, 32'hc16ec1be} /* (11, 9, 20) {real, imag} */,
  {32'hbd9ce600, 32'hbf9f9ea0} /* (11, 9, 19) {real, imag} */,
  {32'h423ed226, 32'h413243e5} /* (11, 9, 18) {real, imag} */,
  {32'h409b86d6, 32'hc2388b2e} /* (11, 9, 17) {real, imag} */,
  {32'hc20ddcc4, 32'h00000000} /* (11, 9, 16) {real, imag} */,
  {32'h409b86d6, 32'h42388b2e} /* (11, 9, 15) {real, imag} */,
  {32'h423ed226, 32'hc13243e5} /* (11, 9, 14) {real, imag} */,
  {32'hbd9ce600, 32'h3f9f9ea0} /* (11, 9, 13) {real, imag} */,
  {32'hc2779c3c, 32'h416ec1be} /* (11, 9, 12) {real, imag} */,
  {32'h4246375a, 32'hc1d90570} /* (11, 9, 11) {real, imag} */,
  {32'h429e5754, 32'hc2a54814} /* (11, 9, 10) {real, imag} */,
  {32'h42bcbf9e, 32'h41c90fa4} /* (11, 9, 9) {real, imag} */,
  {32'hc24db223, 32'h3f3d5ba0} /* (11, 9, 8) {real, imag} */,
  {32'h4227a76c, 32'h41b9c792} /* (11, 9, 7) {real, imag} */,
  {32'hc27fedb1, 32'hc2aa8596} /* (11, 9, 6) {real, imag} */,
  {32'hc2cb68b0, 32'hc32ee31e} /* (11, 9, 5) {real, imag} */,
  {32'h41c023e4, 32'h42d756eb} /* (11, 9, 4) {real, imag} */,
  {32'hc2a89b66, 32'h4334ee74} /* (11, 9, 3) {real, imag} */,
  {32'hc44e1142, 32'hc39a51d4} /* (11, 9, 2) {real, imag} */,
  {32'h44e5fbec, 32'h44856cca} /* (11, 9, 1) {real, imag} */,
  {32'h45270ea7, 32'h00000000} /* (11, 9, 0) {real, imag} */,
  {32'h45288c0e, 32'hc4b82421} /* (11, 8, 31) {real, imag} */,
  {32'hc481fbe8, 32'h43c81375} /* (11, 8, 30) {real, imag} */,
  {32'hc29348f1, 32'hbfad8b20} /* (11, 8, 29) {real, imag} */,
  {32'hc22504ee, 32'h408ea248} /* (11, 8, 28) {real, imag} */,
  {32'hc1f1a7d0, 32'h433289a6} /* (11, 8, 27) {real, imag} */,
  {32'hc1156e08, 32'h42b3c908} /* (11, 8, 26) {real, imag} */,
  {32'h42ddfec6, 32'hc1fda4dc} /* (11, 8, 25) {real, imag} */,
  {32'hc1753754, 32'h423f8ab7} /* (11, 8, 24) {real, imag} */,
  {32'hc2bde8cc, 32'h42bcd9f2} /* (11, 8, 23) {real, imag} */,
  {32'h41e8a05a, 32'h42b5d450} /* (11, 8, 22) {real, imag} */,
  {32'hc2335a38, 32'hc2aae65b} /* (11, 8, 21) {real, imag} */,
  {32'h42c52680, 32'h40126a30} /* (11, 8, 20) {real, imag} */,
  {32'h41c06ded, 32'h42e1c5a5} /* (11, 8, 19) {real, imag} */,
  {32'hc1727b64, 32'h4228170c} /* (11, 8, 18) {real, imag} */,
  {32'hc18100ec, 32'hc1f39bee} /* (11, 8, 17) {real, imag} */,
  {32'h4280a0dc, 32'h00000000} /* (11, 8, 16) {real, imag} */,
  {32'hc18100ec, 32'h41f39bee} /* (11, 8, 15) {real, imag} */,
  {32'hc1727b64, 32'hc228170c} /* (11, 8, 14) {real, imag} */,
  {32'h41c06ded, 32'hc2e1c5a5} /* (11, 8, 13) {real, imag} */,
  {32'h42c52680, 32'hc0126a30} /* (11, 8, 12) {real, imag} */,
  {32'hc2335a38, 32'h42aae65b} /* (11, 8, 11) {real, imag} */,
  {32'h41e8a05a, 32'hc2b5d450} /* (11, 8, 10) {real, imag} */,
  {32'hc2bde8cc, 32'hc2bcd9f2} /* (11, 8, 9) {real, imag} */,
  {32'hc1753754, 32'hc23f8ab7} /* (11, 8, 8) {real, imag} */,
  {32'h42ddfec6, 32'h41fda4dc} /* (11, 8, 7) {real, imag} */,
  {32'hc1156e08, 32'hc2b3c908} /* (11, 8, 6) {real, imag} */,
  {32'hc1f1a7d0, 32'hc33289a6} /* (11, 8, 5) {real, imag} */,
  {32'hc22504ee, 32'hc08ea248} /* (11, 8, 4) {real, imag} */,
  {32'hc29348f1, 32'h3fad8b20} /* (11, 8, 3) {real, imag} */,
  {32'hc481fbe8, 32'hc3c81375} /* (11, 8, 2) {real, imag} */,
  {32'h45288c0e, 32'h44b82421} /* (11, 8, 1) {real, imag} */,
  {32'h455dfc1c, 32'h00000000} /* (11, 8, 0) {real, imag} */,
  {32'h454bb402, 32'hc4e0965c} /* (11, 7, 31) {real, imag} */,
  {32'hc48f0cc0, 32'h44442982} /* (11, 7, 30) {real, imag} */,
  {32'hc3089056, 32'h41886258} /* (11, 7, 29) {real, imag} */,
  {32'hc181219e, 32'hc282199f} /* (11, 7, 28) {real, imag} */,
  {32'hc293228b, 32'h4338830e} /* (11, 7, 27) {real, imag} */,
  {32'h41e9c7e8, 32'hc1dd3980} /* (11, 7, 26) {real, imag} */,
  {32'hc2a2fb27, 32'hc2da1eda} /* (11, 7, 25) {real, imag} */,
  {32'hc2a2a13c, 32'hc1686ff8} /* (11, 7, 24) {real, imag} */,
  {32'hc1093a14, 32'hc2f07473} /* (11, 7, 23) {real, imag} */,
  {32'hc127e314, 32'hc1f0d704} /* (11, 7, 22) {real, imag} */,
  {32'h415b521c, 32'h4180b948} /* (11, 7, 21) {real, imag} */,
  {32'h418f2242, 32'hc1aa66c6} /* (11, 7, 20) {real, imag} */,
  {32'h421a30e5, 32'hc2a27291} /* (11, 7, 19) {real, imag} */,
  {32'hbec44f40, 32'hc19c5e66} /* (11, 7, 18) {real, imag} */,
  {32'h416174c3, 32'h420ad10c} /* (11, 7, 17) {real, imag} */,
  {32'hc2df2c3c, 32'h00000000} /* (11, 7, 16) {real, imag} */,
  {32'h416174c3, 32'hc20ad10c} /* (11, 7, 15) {real, imag} */,
  {32'hbec44f40, 32'h419c5e66} /* (11, 7, 14) {real, imag} */,
  {32'h421a30e5, 32'h42a27291} /* (11, 7, 13) {real, imag} */,
  {32'h418f2242, 32'h41aa66c6} /* (11, 7, 12) {real, imag} */,
  {32'h415b521c, 32'hc180b948} /* (11, 7, 11) {real, imag} */,
  {32'hc127e314, 32'h41f0d704} /* (11, 7, 10) {real, imag} */,
  {32'hc1093a14, 32'h42f07473} /* (11, 7, 9) {real, imag} */,
  {32'hc2a2a13c, 32'h41686ff8} /* (11, 7, 8) {real, imag} */,
  {32'hc2a2fb27, 32'h42da1eda} /* (11, 7, 7) {real, imag} */,
  {32'h41e9c7e8, 32'h41dd3980} /* (11, 7, 6) {real, imag} */,
  {32'hc293228b, 32'hc338830e} /* (11, 7, 5) {real, imag} */,
  {32'hc181219e, 32'h4282199f} /* (11, 7, 4) {real, imag} */,
  {32'hc3089056, 32'hc1886258} /* (11, 7, 3) {real, imag} */,
  {32'hc48f0cc0, 32'hc4442982} /* (11, 7, 2) {real, imag} */,
  {32'h454bb402, 32'h44e0965c} /* (11, 7, 1) {real, imag} */,
  {32'h4587d105, 32'h00000000} /* (11, 7, 0) {real, imag} */,
  {32'h4563f9fe, 32'hc50ded8b} /* (11, 6, 31) {real, imag} */,
  {32'hc471d296, 32'h44626d2c} /* (11, 6, 30) {real, imag} */,
  {32'hc301cf78, 32'hc27634d6} /* (11, 6, 29) {real, imag} */,
  {32'h4304d311, 32'hc1d17fca} /* (11, 6, 28) {real, imag} */,
  {32'hc17bb5f8, 32'h43ac66ac} /* (11, 6, 27) {real, imag} */,
  {32'hc1212dfc, 32'hc2300c18} /* (11, 6, 26) {real, imag} */,
  {32'hc23286b8, 32'hc267c09d} /* (11, 6, 25) {real, imag} */,
  {32'h4261b9ae, 32'hc21a1fcc} /* (11, 6, 24) {real, imag} */,
  {32'h42082afc, 32'h4190fc78} /* (11, 6, 23) {real, imag} */,
  {32'hc176413c, 32'h42e79725} /* (11, 6, 22) {real, imag} */,
  {32'hc296f14f, 32'h421040b0} /* (11, 6, 21) {real, imag} */,
  {32'h420c0a8a, 32'hc02200f4} /* (11, 6, 20) {real, imag} */,
  {32'hc2b48d0e, 32'hc1a2d488} /* (11, 6, 19) {real, imag} */,
  {32'hc2c9a4f1, 32'h42ab30b0} /* (11, 6, 18) {real, imag} */,
  {32'h4300da10, 32'hc2778d34} /* (11, 6, 17) {real, imag} */,
  {32'hc12db9c7, 32'h00000000} /* (11, 6, 16) {real, imag} */,
  {32'h4300da10, 32'h42778d34} /* (11, 6, 15) {real, imag} */,
  {32'hc2c9a4f1, 32'hc2ab30b0} /* (11, 6, 14) {real, imag} */,
  {32'hc2b48d0e, 32'h41a2d488} /* (11, 6, 13) {real, imag} */,
  {32'h420c0a8a, 32'h402200f4} /* (11, 6, 12) {real, imag} */,
  {32'hc296f14f, 32'hc21040b0} /* (11, 6, 11) {real, imag} */,
  {32'hc176413c, 32'hc2e79725} /* (11, 6, 10) {real, imag} */,
  {32'h42082afc, 32'hc190fc78} /* (11, 6, 9) {real, imag} */,
  {32'h4261b9ae, 32'h421a1fcc} /* (11, 6, 8) {real, imag} */,
  {32'hc23286b8, 32'h4267c09d} /* (11, 6, 7) {real, imag} */,
  {32'hc1212dfc, 32'h42300c18} /* (11, 6, 6) {real, imag} */,
  {32'hc17bb5f8, 32'hc3ac66ac} /* (11, 6, 5) {real, imag} */,
  {32'h4304d311, 32'h41d17fca} /* (11, 6, 4) {real, imag} */,
  {32'hc301cf78, 32'h427634d6} /* (11, 6, 3) {real, imag} */,
  {32'hc471d296, 32'hc4626d2c} /* (11, 6, 2) {real, imag} */,
  {32'h4563f9fe, 32'h450ded8b} /* (11, 6, 1) {real, imag} */,
  {32'h45939a96, 32'h00000000} /* (11, 6, 0) {real, imag} */,
  {32'h4558882e, 32'hc544569a} /* (11, 5, 31) {real, imag} */,
  {32'hc3bdb656, 32'h448370ea} /* (11, 5, 30) {real, imag} */,
  {32'hc28d4df4, 32'hc098c720} /* (11, 5, 29) {real, imag} */,
  {32'hc188a920, 32'h43931310} /* (11, 5, 28) {real, imag} */,
  {32'hc3000df8, 32'h432f33e2} /* (11, 5, 27) {real, imag} */,
  {32'hc2ff891e, 32'h42e2a8c0} /* (11, 5, 26) {real, imag} */,
  {32'h42bbbcff, 32'hc30ca2c0} /* (11, 5, 25) {real, imag} */,
  {32'hc2196676, 32'hc2322e75} /* (11, 5, 24) {real, imag} */,
  {32'hc2dc2b7c, 32'h4300d962} /* (11, 5, 23) {real, imag} */,
  {32'h42364b54, 32'h41b4198c} /* (11, 5, 22) {real, imag} */,
  {32'hc2441eba, 32'h4301c14e} /* (11, 5, 21) {real, imag} */,
  {32'h42272bd8, 32'hc292a601} /* (11, 5, 20) {real, imag} */,
  {32'h42a46517, 32'h423da068} /* (11, 5, 19) {real, imag} */,
  {32'hc2941577, 32'hc10ae22c} /* (11, 5, 18) {real, imag} */,
  {32'hc248d605, 32'hc1fbb98c} /* (11, 5, 17) {real, imag} */,
  {32'hc28c5ca6, 32'h00000000} /* (11, 5, 16) {real, imag} */,
  {32'hc248d605, 32'h41fbb98c} /* (11, 5, 15) {real, imag} */,
  {32'hc2941577, 32'h410ae22c} /* (11, 5, 14) {real, imag} */,
  {32'h42a46517, 32'hc23da068} /* (11, 5, 13) {real, imag} */,
  {32'h42272bd8, 32'h4292a601} /* (11, 5, 12) {real, imag} */,
  {32'hc2441eba, 32'hc301c14e} /* (11, 5, 11) {real, imag} */,
  {32'h42364b54, 32'hc1b4198c} /* (11, 5, 10) {real, imag} */,
  {32'hc2dc2b7c, 32'hc300d962} /* (11, 5, 9) {real, imag} */,
  {32'hc2196676, 32'h42322e75} /* (11, 5, 8) {real, imag} */,
  {32'h42bbbcff, 32'h430ca2c0} /* (11, 5, 7) {real, imag} */,
  {32'hc2ff891e, 32'hc2e2a8c0} /* (11, 5, 6) {real, imag} */,
  {32'hc3000df8, 32'hc32f33e2} /* (11, 5, 5) {real, imag} */,
  {32'hc188a920, 32'hc3931310} /* (11, 5, 4) {real, imag} */,
  {32'hc28d4df4, 32'h4098c720} /* (11, 5, 3) {real, imag} */,
  {32'hc3bdb656, 32'hc48370ea} /* (11, 5, 2) {real, imag} */,
  {32'h4558882e, 32'h4544569a} /* (11, 5, 1) {real, imag} */,
  {32'h45a29b4a, 32'h00000000} /* (11, 5, 0) {real, imag} */,
  {32'h453ce750, 32'hc56c6448} /* (11, 4, 31) {real, imag} */,
  {32'h430e30b8, 32'h44a68d34} /* (11, 4, 30) {real, imag} */,
  {32'hc2a20c4d, 32'h41fb2cf8} /* (11, 4, 29) {real, imag} */,
  {32'hc313fca8, 32'h435b073a} /* (11, 4, 28) {real, imag} */,
  {32'hc3610d2a, 32'hc2d60b20} /* (11, 4, 27) {real, imag} */,
  {32'h41861a18, 32'h425b9080} /* (11, 4, 26) {real, imag} */,
  {32'hc28e103a, 32'hc264546d} /* (11, 4, 25) {real, imag} */,
  {32'hc241b4f5, 32'h431f7878} /* (11, 4, 24) {real, imag} */,
  {32'hc22200b6, 32'hc26f0550} /* (11, 4, 23) {real, imag} */,
  {32'h4316f171, 32'h41a2049c} /* (11, 4, 22) {real, imag} */,
  {32'hc264442c, 32'hc193aa9d} /* (11, 4, 21) {real, imag} */,
  {32'hc2473ce8, 32'h428f3e81} /* (11, 4, 20) {real, imag} */,
  {32'h427f1afb, 32'h413374aa} /* (11, 4, 19) {real, imag} */,
  {32'h4293dfe6, 32'h42413840} /* (11, 4, 18) {real, imag} */,
  {32'hc2957354, 32'hc1eec611} /* (11, 4, 17) {real, imag} */,
  {32'hc05b7140, 32'h00000000} /* (11, 4, 16) {real, imag} */,
  {32'hc2957354, 32'h41eec611} /* (11, 4, 15) {real, imag} */,
  {32'h4293dfe6, 32'hc2413840} /* (11, 4, 14) {real, imag} */,
  {32'h427f1afb, 32'hc13374aa} /* (11, 4, 13) {real, imag} */,
  {32'hc2473ce8, 32'hc28f3e81} /* (11, 4, 12) {real, imag} */,
  {32'hc264442c, 32'h4193aa9d} /* (11, 4, 11) {real, imag} */,
  {32'h4316f171, 32'hc1a2049c} /* (11, 4, 10) {real, imag} */,
  {32'hc22200b6, 32'h426f0550} /* (11, 4, 9) {real, imag} */,
  {32'hc241b4f5, 32'hc31f7878} /* (11, 4, 8) {real, imag} */,
  {32'hc28e103a, 32'h4264546d} /* (11, 4, 7) {real, imag} */,
  {32'h41861a18, 32'hc25b9080} /* (11, 4, 6) {real, imag} */,
  {32'hc3610d2a, 32'h42d60b20} /* (11, 4, 5) {real, imag} */,
  {32'hc313fca8, 32'hc35b073a} /* (11, 4, 4) {real, imag} */,
  {32'hc2a20c4d, 32'hc1fb2cf8} /* (11, 4, 3) {real, imag} */,
  {32'h430e30b8, 32'hc4a68d34} /* (11, 4, 2) {real, imag} */,
  {32'h453ce750, 32'h456c6448} /* (11, 4, 1) {real, imag} */,
  {32'h45b0555a, 32'h00000000} /* (11, 4, 0) {real, imag} */,
  {32'h4546af41, 32'hc57ec301} /* (11, 3, 31) {real, imag} */,
  {32'h437a0814, 32'h448ef4be} /* (11, 3, 30) {real, imag} */,
  {32'hc2c23cc6, 32'hc234ddca} /* (11, 3, 29) {real, imag} */,
  {32'hc32a6e72, 32'h436ab9fe} /* (11, 3, 28) {real, imag} */,
  {32'hc3758d2e, 32'hc2b5d2ff} /* (11, 3, 27) {real, imag} */,
  {32'hc266ed88, 32'h42852599} /* (11, 3, 26) {real, imag} */,
  {32'hc20d0264, 32'h413dcce8} /* (11, 3, 25) {real, imag} */,
  {32'h41fca5ee, 32'h42cf4001} /* (11, 3, 24) {real, imag} */,
  {32'h422798e4, 32'h428a4f96} /* (11, 3, 23) {real, imag} */,
  {32'h4218feb8, 32'h423f900e} /* (11, 3, 22) {real, imag} */,
  {32'hc2a1cfcf, 32'hc215df2a} /* (11, 3, 21) {real, imag} */,
  {32'hc11fb56b, 32'h41d6c49e} /* (11, 3, 20) {real, imag} */,
  {32'hc222c0f8, 32'hc3152d12} /* (11, 3, 19) {real, imag} */,
  {32'h42b5dff0, 32'hc1c002f4} /* (11, 3, 18) {real, imag} */,
  {32'hc22edfb6, 32'h4100c9e2} /* (11, 3, 17) {real, imag} */,
  {32'hc0ce491c, 32'h00000000} /* (11, 3, 16) {real, imag} */,
  {32'hc22edfb6, 32'hc100c9e2} /* (11, 3, 15) {real, imag} */,
  {32'h42b5dff0, 32'h41c002f4} /* (11, 3, 14) {real, imag} */,
  {32'hc222c0f8, 32'h43152d12} /* (11, 3, 13) {real, imag} */,
  {32'hc11fb56b, 32'hc1d6c49e} /* (11, 3, 12) {real, imag} */,
  {32'hc2a1cfcf, 32'h4215df2a} /* (11, 3, 11) {real, imag} */,
  {32'h4218feb8, 32'hc23f900e} /* (11, 3, 10) {real, imag} */,
  {32'h422798e4, 32'hc28a4f96} /* (11, 3, 9) {real, imag} */,
  {32'h41fca5ee, 32'hc2cf4001} /* (11, 3, 8) {real, imag} */,
  {32'hc20d0264, 32'hc13dcce8} /* (11, 3, 7) {real, imag} */,
  {32'hc266ed88, 32'hc2852599} /* (11, 3, 6) {real, imag} */,
  {32'hc3758d2e, 32'h42b5d2ff} /* (11, 3, 5) {real, imag} */,
  {32'hc32a6e72, 32'hc36ab9fe} /* (11, 3, 4) {real, imag} */,
  {32'hc2c23cc6, 32'h4234ddca} /* (11, 3, 3) {real, imag} */,
  {32'h437a0814, 32'hc48ef4be} /* (11, 3, 2) {real, imag} */,
  {32'h4546af41, 32'h457ec301} /* (11, 3, 1) {real, imag} */,
  {32'h45ae2263, 32'h00000000} /* (11, 3, 0) {real, imag} */,
  {32'h454e644a, 32'hc57ce094} /* (11, 2, 31) {real, imag} */,
  {32'h4381981a, 32'h448e95dd} /* (11, 2, 30) {real, imag} */,
  {32'hc2331baa, 32'hc0d80c58} /* (11, 2, 29) {real, imag} */,
  {32'hc34f1ba4, 32'h43ac5bdc} /* (11, 2, 28) {real, imag} */,
  {32'hc380a36c, 32'hc2890c33} /* (11, 2, 27) {real, imag} */,
  {32'hc31113c6, 32'h41828d68} /* (11, 2, 26) {real, imag} */,
  {32'h415ea0dc, 32'hc0eaa828} /* (11, 2, 25) {real, imag} */,
  {32'h4311dd34, 32'h415a57e8} /* (11, 2, 24) {real, imag} */,
  {32'hbf960e60, 32'hc0b24c88} /* (11, 2, 23) {real, imag} */,
  {32'hc28d2aa8, 32'h42acfc09} /* (11, 2, 22) {real, imag} */,
  {32'hc1f9f58a, 32'hc2560cd0} /* (11, 2, 21) {real, imag} */,
  {32'hc2e8b59a, 32'hc233280a} /* (11, 2, 20) {real, imag} */,
  {32'hc25fb0fa, 32'hc262e5a7} /* (11, 2, 19) {real, imag} */,
  {32'h42566bcb, 32'h41f04e52} /* (11, 2, 18) {real, imag} */,
  {32'h41ea59b5, 32'hc1b1732b} /* (11, 2, 17) {real, imag} */,
  {32'hc2017f78, 32'h00000000} /* (11, 2, 16) {real, imag} */,
  {32'h41ea59b5, 32'h41b1732b} /* (11, 2, 15) {real, imag} */,
  {32'h42566bcb, 32'hc1f04e52} /* (11, 2, 14) {real, imag} */,
  {32'hc25fb0fa, 32'h4262e5a7} /* (11, 2, 13) {real, imag} */,
  {32'hc2e8b59a, 32'h4233280a} /* (11, 2, 12) {real, imag} */,
  {32'hc1f9f58a, 32'h42560cd0} /* (11, 2, 11) {real, imag} */,
  {32'hc28d2aa8, 32'hc2acfc09} /* (11, 2, 10) {real, imag} */,
  {32'hbf960e60, 32'h40b24c88} /* (11, 2, 9) {real, imag} */,
  {32'h4311dd34, 32'hc15a57e8} /* (11, 2, 8) {real, imag} */,
  {32'h415ea0dc, 32'h40eaa828} /* (11, 2, 7) {real, imag} */,
  {32'hc31113c6, 32'hc1828d68} /* (11, 2, 6) {real, imag} */,
  {32'hc380a36c, 32'h42890c33} /* (11, 2, 5) {real, imag} */,
  {32'hc34f1ba4, 32'hc3ac5bdc} /* (11, 2, 4) {real, imag} */,
  {32'hc2331baa, 32'h40d80c58} /* (11, 2, 3) {real, imag} */,
  {32'h4381981a, 32'hc48e95dd} /* (11, 2, 2) {real, imag} */,
  {32'h454e644a, 32'h457ce094} /* (11, 2, 1) {real, imag} */,
  {32'h45acc3c1, 32'h00000000} /* (11, 2, 0) {real, imag} */,
  {32'h4556c645, 32'hc56b2684} /* (11, 1, 31) {real, imag} */,
  {32'h41f975a0, 32'h44658441} /* (11, 1, 30) {real, imag} */,
  {32'hc2e87718, 32'hc27aec52} /* (11, 1, 29) {real, imag} */,
  {32'hc326201c, 32'h43889cd6} /* (11, 1, 28) {real, imag} */,
  {32'hc328681a, 32'hc2a44c48} /* (11, 1, 27) {real, imag} */,
  {32'hc239430e, 32'hbfca2b60} /* (11, 1, 26) {real, imag} */,
  {32'h42fb4a52, 32'h428a2af4} /* (11, 1, 25) {real, imag} */,
  {32'h42a6922b, 32'h4213e642} /* (11, 1, 24) {real, imag} */,
  {32'hc27e5b56, 32'h40a1bbe4} /* (11, 1, 23) {real, imag} */,
  {32'hc24b4343, 32'h42c1ce9e} /* (11, 1, 22) {real, imag} */,
  {32'h41e414f8, 32'h419af38e} /* (11, 1, 21) {real, imag} */,
  {32'h4286ac02, 32'hc0aa04ec} /* (11, 1, 20) {real, imag} */,
  {32'hc282c902, 32'h428e390d} /* (11, 1, 19) {real, imag} */,
  {32'h42296b4d, 32'hc1d53664} /* (11, 1, 18) {real, imag} */,
  {32'hc215fa2d, 32'h41ce4715} /* (11, 1, 17) {real, imag} */,
  {32'h41eb74fa, 32'h00000000} /* (11, 1, 16) {real, imag} */,
  {32'hc215fa2d, 32'hc1ce4715} /* (11, 1, 15) {real, imag} */,
  {32'h42296b4d, 32'h41d53664} /* (11, 1, 14) {real, imag} */,
  {32'hc282c902, 32'hc28e390d} /* (11, 1, 13) {real, imag} */,
  {32'h4286ac02, 32'h40aa04ec} /* (11, 1, 12) {real, imag} */,
  {32'h41e414f8, 32'hc19af38e} /* (11, 1, 11) {real, imag} */,
  {32'hc24b4343, 32'hc2c1ce9e} /* (11, 1, 10) {real, imag} */,
  {32'hc27e5b56, 32'hc0a1bbe4} /* (11, 1, 9) {real, imag} */,
  {32'h42a6922b, 32'hc213e642} /* (11, 1, 8) {real, imag} */,
  {32'h42fb4a52, 32'hc28a2af4} /* (11, 1, 7) {real, imag} */,
  {32'hc239430e, 32'h3fca2b60} /* (11, 1, 6) {real, imag} */,
  {32'hc328681a, 32'h42a44c48} /* (11, 1, 5) {real, imag} */,
  {32'hc326201c, 32'hc3889cd6} /* (11, 1, 4) {real, imag} */,
  {32'hc2e87718, 32'h427aec52} /* (11, 1, 3) {real, imag} */,
  {32'h41f975a0, 32'hc4658441} /* (11, 1, 2) {real, imag} */,
  {32'h4556c645, 32'h456b2684} /* (11, 1, 1) {real, imag} */,
  {32'h45aff029, 32'h00000000} /* (11, 1, 0) {real, imag} */,
  {32'h455f585d, 32'hc53ec240} /* (11, 0, 31) {real, imag} */,
  {32'hc37ae2c8, 32'h44357374} /* (11, 0, 30) {real, imag} */,
  {32'hc2c71d06, 32'h40eb32a8} /* (11, 0, 29) {real, imag} */,
  {32'hc2408f62, 32'h43844a58} /* (11, 0, 28) {real, imag} */,
  {32'hc30fc678, 32'hc2714990} /* (11, 0, 27) {real, imag} */,
  {32'h412faa1c, 32'h4292fc0b} /* (11, 0, 26) {real, imag} */,
  {32'h42ae3f6c, 32'h42269cec} /* (11, 0, 25) {real, imag} */,
  {32'h419b300b, 32'h40441fc0} /* (11, 0, 24) {real, imag} */,
  {32'hc2847834, 32'h4176d9cc} /* (11, 0, 23) {real, imag} */,
  {32'h4020a3c0, 32'hc2176552} /* (11, 0, 22) {real, imag} */,
  {32'hc23a1a22, 32'h4214e170} /* (11, 0, 21) {real, imag} */,
  {32'h4245405e, 32'h41cf4230} /* (11, 0, 20) {real, imag} */,
  {32'hc131e72c, 32'h40745b00} /* (11, 0, 19) {real, imag} */,
  {32'h41987108, 32'hc06b7910} /* (11, 0, 18) {real, imag} */,
  {32'hc0141d48, 32'h40b4d244} /* (11, 0, 17) {real, imag} */,
  {32'hc2a3a182, 32'h00000000} /* (11, 0, 16) {real, imag} */,
  {32'hc0141d48, 32'hc0b4d244} /* (11, 0, 15) {real, imag} */,
  {32'h41987108, 32'h406b7910} /* (11, 0, 14) {real, imag} */,
  {32'hc131e72c, 32'hc0745b00} /* (11, 0, 13) {real, imag} */,
  {32'h4245405e, 32'hc1cf4230} /* (11, 0, 12) {real, imag} */,
  {32'hc23a1a22, 32'hc214e170} /* (11, 0, 11) {real, imag} */,
  {32'h4020a3c0, 32'h42176552} /* (11, 0, 10) {real, imag} */,
  {32'hc2847834, 32'hc176d9cc} /* (11, 0, 9) {real, imag} */,
  {32'h419b300b, 32'hc0441fc0} /* (11, 0, 8) {real, imag} */,
  {32'h42ae3f6c, 32'hc2269cec} /* (11, 0, 7) {real, imag} */,
  {32'h412faa1c, 32'hc292fc0b} /* (11, 0, 6) {real, imag} */,
  {32'hc30fc678, 32'h42714990} /* (11, 0, 5) {real, imag} */,
  {32'hc2408f62, 32'hc3844a58} /* (11, 0, 4) {real, imag} */,
  {32'hc2c71d06, 32'hc0eb32a8} /* (11, 0, 3) {real, imag} */,
  {32'hc37ae2c8, 32'hc4357374} /* (11, 0, 2) {real, imag} */,
  {32'h455f585d, 32'h453ec240} /* (11, 0, 1) {real, imag} */,
  {32'h45ac3538, 32'h00000000} /* (11, 0, 0) {real, imag} */,
  {32'h4580f03b, 32'hc518cf90} /* (10, 31, 31) {real, imag} */,
  {32'hc454b627, 32'h44469b0e} /* (10, 31, 30) {real, imag} */,
  {32'hc0346ea0, 32'hc22e20ef} /* (10, 31, 29) {real, imag} */,
  {32'h4310d49a, 32'h420c2e20} /* (10, 31, 28) {real, imag} */,
  {32'hc301bdfc, 32'hc1b267ac} /* (10, 31, 27) {real, imag} */,
  {32'h41ef7eeb, 32'h43055efe} /* (10, 31, 26) {real, imag} */,
  {32'h424ee255, 32'h4136b9e8} /* (10, 31, 25) {real, imag} */,
  {32'hc22713be, 32'h427fe6a7} /* (10, 31, 24) {real, imag} */,
  {32'h429c96bc, 32'hc10f7858} /* (10, 31, 23) {real, imag} */,
  {32'hc1934bfc, 32'h41a8e942} /* (10, 31, 22) {real, imag} */,
  {32'h419df37e, 32'h41e166aa} /* (10, 31, 21) {real, imag} */,
  {32'h41194538, 32'h431091d6} /* (10, 31, 20) {real, imag} */,
  {32'hc1bd73f3, 32'hc0eb0974} /* (10, 31, 19) {real, imag} */,
  {32'hc138286c, 32'hbffa8a60} /* (10, 31, 18) {real, imag} */,
  {32'hc0588d80, 32'hc233fb30} /* (10, 31, 17) {real, imag} */,
  {32'hc130c1d8, 32'h00000000} /* (10, 31, 16) {real, imag} */,
  {32'hc0588d80, 32'h4233fb30} /* (10, 31, 15) {real, imag} */,
  {32'hc138286c, 32'h3ffa8a60} /* (10, 31, 14) {real, imag} */,
  {32'hc1bd73f3, 32'h40eb0974} /* (10, 31, 13) {real, imag} */,
  {32'h41194538, 32'hc31091d6} /* (10, 31, 12) {real, imag} */,
  {32'h419df37e, 32'hc1e166aa} /* (10, 31, 11) {real, imag} */,
  {32'hc1934bfc, 32'hc1a8e942} /* (10, 31, 10) {real, imag} */,
  {32'h429c96bc, 32'h410f7858} /* (10, 31, 9) {real, imag} */,
  {32'hc22713be, 32'hc27fe6a7} /* (10, 31, 8) {real, imag} */,
  {32'h424ee255, 32'hc136b9e8} /* (10, 31, 7) {real, imag} */,
  {32'h41ef7eeb, 32'hc3055efe} /* (10, 31, 6) {real, imag} */,
  {32'hc301bdfc, 32'h41b267ac} /* (10, 31, 5) {real, imag} */,
  {32'h4310d49a, 32'hc20c2e20} /* (10, 31, 4) {real, imag} */,
  {32'hc0346ea0, 32'h422e20ef} /* (10, 31, 3) {real, imag} */,
  {32'hc454b627, 32'hc4469b0e} /* (10, 31, 2) {real, imag} */,
  {32'h4580f03b, 32'h4518cf90} /* (10, 31, 1) {real, imag} */,
  {32'h45b1c50f, 32'h00000000} /* (10, 31, 0) {real, imag} */,
  {32'h4593f067, 32'hc4ec31ca} /* (10, 30, 31) {real, imag} */,
  {32'hc49828da, 32'h442d9d26} /* (10, 30, 30) {real, imag} */,
  {32'hc00abc20, 32'hc30dc6d4} /* (10, 30, 29) {real, imag} */,
  {32'h43463534, 32'h40d79560} /* (10, 30, 28) {real, imag} */,
  {32'hc3699034, 32'h423f2b7d} /* (10, 30, 27) {real, imag} */,
  {32'hc2585fb7, 32'h41b5fb28} /* (10, 30, 26) {real, imag} */,
  {32'h41439e72, 32'hc1402a00} /* (10, 30, 25) {real, imag} */,
  {32'hc0eb7748, 32'h4245833d} /* (10, 30, 24) {real, imag} */,
  {32'h421ce365, 32'h4223800f} /* (10, 30, 23) {real, imag} */,
  {32'hc3115f7e, 32'h41918efc} /* (10, 30, 22) {real, imag} */,
  {32'hc2a027e9, 32'hc2796a84} /* (10, 30, 21) {real, imag} */,
  {32'hc1f0e658, 32'h428162d9} /* (10, 30, 20) {real, imag} */,
  {32'hc0bf6746, 32'h41fda1ac} /* (10, 30, 19) {real, imag} */,
  {32'hc295d5b4, 32'h41b60816} /* (10, 30, 18) {real, imag} */,
  {32'h426b0f87, 32'h4145dcc9} /* (10, 30, 17) {real, imag} */,
  {32'h417ca7e4, 32'h00000000} /* (10, 30, 16) {real, imag} */,
  {32'h426b0f87, 32'hc145dcc9} /* (10, 30, 15) {real, imag} */,
  {32'hc295d5b4, 32'hc1b60816} /* (10, 30, 14) {real, imag} */,
  {32'hc0bf6746, 32'hc1fda1ac} /* (10, 30, 13) {real, imag} */,
  {32'hc1f0e658, 32'hc28162d9} /* (10, 30, 12) {real, imag} */,
  {32'hc2a027e9, 32'h42796a84} /* (10, 30, 11) {real, imag} */,
  {32'hc3115f7e, 32'hc1918efc} /* (10, 30, 10) {real, imag} */,
  {32'h421ce365, 32'hc223800f} /* (10, 30, 9) {real, imag} */,
  {32'hc0eb7748, 32'hc245833d} /* (10, 30, 8) {real, imag} */,
  {32'h41439e72, 32'h41402a00} /* (10, 30, 7) {real, imag} */,
  {32'hc2585fb7, 32'hc1b5fb28} /* (10, 30, 6) {real, imag} */,
  {32'hc3699034, 32'hc23f2b7d} /* (10, 30, 5) {real, imag} */,
  {32'h43463534, 32'hc0d79560} /* (10, 30, 4) {real, imag} */,
  {32'hc00abc20, 32'h430dc6d4} /* (10, 30, 3) {real, imag} */,
  {32'hc49828da, 32'hc42d9d26} /* (10, 30, 2) {real, imag} */,
  {32'h4593f067, 32'h44ec31ca} /* (10, 30, 1) {real, imag} */,
  {32'h45b7c5f9, 32'h00000000} /* (10, 30, 0) {real, imag} */,
  {32'h459dd546, 32'hc4b316ef} /* (10, 29, 31) {real, imag} */,
  {32'hc4afa18c, 32'h43fe0bc5} /* (10, 29, 30) {real, imag} */,
  {32'hc1543ef8, 32'hc1456024} /* (10, 29, 29) {real, imag} */,
  {32'h434737f2, 32'hc2146870} /* (10, 29, 28) {real, imag} */,
  {32'hc3265b1e, 32'h42978710} /* (10, 29, 27) {real, imag} */,
  {32'hc0d8bb88, 32'hc289dd90} /* (10, 29, 26) {real, imag} */,
  {32'hc0514c84, 32'hc30a94c4} /* (10, 29, 25) {real, imag} */,
  {32'hc236b42c, 32'h421856bc} /* (10, 29, 24) {real, imag} */,
  {32'hc07afc9c, 32'hc1a1d2f8} /* (10, 29, 23) {real, imag} */,
  {32'h426f0a6b, 32'h42d0241e} /* (10, 29, 22) {real, imag} */,
  {32'hc25b2780, 32'h424721c4} /* (10, 29, 21) {real, imag} */,
  {32'h41e7ee84, 32'hc1c0411a} /* (10, 29, 20) {real, imag} */,
  {32'hc0a08860, 32'hc1477738} /* (10, 29, 19) {real, imag} */,
  {32'hc1401d2c, 32'h42dde944} /* (10, 29, 18) {real, imag} */,
  {32'hc1a63c70, 32'hc1c9f0da} /* (10, 29, 17) {real, imag} */,
  {32'h41a93b74, 32'h00000000} /* (10, 29, 16) {real, imag} */,
  {32'hc1a63c70, 32'h41c9f0da} /* (10, 29, 15) {real, imag} */,
  {32'hc1401d2c, 32'hc2dde944} /* (10, 29, 14) {real, imag} */,
  {32'hc0a08860, 32'h41477738} /* (10, 29, 13) {real, imag} */,
  {32'h41e7ee84, 32'h41c0411a} /* (10, 29, 12) {real, imag} */,
  {32'hc25b2780, 32'hc24721c4} /* (10, 29, 11) {real, imag} */,
  {32'h426f0a6b, 32'hc2d0241e} /* (10, 29, 10) {real, imag} */,
  {32'hc07afc9c, 32'h41a1d2f8} /* (10, 29, 9) {real, imag} */,
  {32'hc236b42c, 32'hc21856bc} /* (10, 29, 8) {real, imag} */,
  {32'hc0514c84, 32'h430a94c4} /* (10, 29, 7) {real, imag} */,
  {32'hc0d8bb88, 32'h4289dd90} /* (10, 29, 6) {real, imag} */,
  {32'hc3265b1e, 32'hc2978710} /* (10, 29, 5) {real, imag} */,
  {32'h434737f2, 32'h42146870} /* (10, 29, 4) {real, imag} */,
  {32'hc1543ef8, 32'h41456024} /* (10, 29, 3) {real, imag} */,
  {32'hc4afa18c, 32'hc3fe0bc5} /* (10, 29, 2) {real, imag} */,
  {32'h459dd546, 32'h44b316ef} /* (10, 29, 1) {real, imag} */,
  {32'h45b8a1ca, 32'h00000000} /* (10, 29, 0) {real, imag} */,
  {32'h45a6b1b6, 32'hc496c8a2} /* (10, 28, 31) {real, imag} */,
  {32'hc4cf4642, 32'h44027b76} /* (10, 28, 30) {real, imag} */,
  {32'hc0d9e120, 32'h42f028e1} /* (10, 28, 29) {real, imag} */,
  {32'h4320701d, 32'hc2923742} /* (10, 28, 28) {real, imag} */,
  {32'hc30686a2, 32'hc2212966} /* (10, 28, 27) {real, imag} */,
  {32'h42310954, 32'h4187c5c2} /* (10, 28, 26) {real, imag} */,
  {32'h42aca3a8, 32'hc1d387f8} /* (10, 28, 25) {real, imag} */,
  {32'hc1a6013b, 32'h42547f80} /* (10, 28, 24) {real, imag} */,
  {32'h40a22588, 32'hc294bae0} /* (10, 28, 23) {real, imag} */,
  {32'h41c8781a, 32'h430204d1} /* (10, 28, 22) {real, imag} */,
  {32'hc2525054, 32'h428e14bc} /* (10, 28, 21) {real, imag} */,
  {32'hc1f95b86, 32'h42aa6660} /* (10, 28, 20) {real, imag} */,
  {32'hc27f819e, 32'hc230204e} /* (10, 28, 19) {real, imag} */,
  {32'hc24e1f12, 32'hc1d2cb7d} /* (10, 28, 18) {real, imag} */,
  {32'h41129772, 32'h42a56e0a} /* (10, 28, 17) {real, imag} */,
  {32'hbf860e8c, 32'h00000000} /* (10, 28, 16) {real, imag} */,
  {32'h41129772, 32'hc2a56e0a} /* (10, 28, 15) {real, imag} */,
  {32'hc24e1f12, 32'h41d2cb7d} /* (10, 28, 14) {real, imag} */,
  {32'hc27f819e, 32'h4230204e} /* (10, 28, 13) {real, imag} */,
  {32'hc1f95b86, 32'hc2aa6660} /* (10, 28, 12) {real, imag} */,
  {32'hc2525054, 32'hc28e14bc} /* (10, 28, 11) {real, imag} */,
  {32'h41c8781a, 32'hc30204d1} /* (10, 28, 10) {real, imag} */,
  {32'h40a22588, 32'h4294bae0} /* (10, 28, 9) {real, imag} */,
  {32'hc1a6013b, 32'hc2547f80} /* (10, 28, 8) {real, imag} */,
  {32'h42aca3a8, 32'h41d387f8} /* (10, 28, 7) {real, imag} */,
  {32'h42310954, 32'hc187c5c2} /* (10, 28, 6) {real, imag} */,
  {32'hc30686a2, 32'h42212966} /* (10, 28, 5) {real, imag} */,
  {32'h4320701d, 32'h42923742} /* (10, 28, 4) {real, imag} */,
  {32'hc0d9e120, 32'hc2f028e1} /* (10, 28, 3) {real, imag} */,
  {32'hc4cf4642, 32'hc4027b76} /* (10, 28, 2) {real, imag} */,
  {32'h45a6b1b6, 32'h4496c8a2} /* (10, 28, 1) {real, imag} */,
  {32'h45b628e2, 32'h00000000} /* (10, 28, 0) {real, imag} */,
  {32'h45aef8f8, 32'hc48aca0f} /* (10, 27, 31) {real, imag} */,
  {32'hc4ec8f80, 32'h439e8ed7} /* (10, 27, 30) {real, imag} */,
  {32'hc21e0849, 32'h4319e569} /* (10, 27, 29) {real, imag} */,
  {32'h42c3923a, 32'hc2d8ce28} /* (10, 27, 28) {real, imag} */,
  {32'hc3165064, 32'hc190605c} /* (10, 27, 27) {real, imag} */,
  {32'h40afeb08, 32'h4181215d} /* (10, 27, 26) {real, imag} */,
  {32'h4334948d, 32'hc2a244dd} /* (10, 27, 25) {real, imag} */,
  {32'hc155a0d0, 32'h42825c40} /* (10, 27, 24) {real, imag} */,
  {32'hc29cb432, 32'h42ebbdfe} /* (10, 27, 23) {real, imag} */,
  {32'h41c44317, 32'h423ab8b9} /* (10, 27, 22) {real, imag} */,
  {32'h42a2a73e, 32'h42eed5b0} /* (10, 27, 21) {real, imag} */,
  {32'h412e6489, 32'hc282bd20} /* (10, 27, 20) {real, imag} */,
  {32'h426f91b5, 32'hc2edab30} /* (10, 27, 19) {real, imag} */,
  {32'h40c646e0, 32'hc298eb06} /* (10, 27, 18) {real, imag} */,
  {32'hc2250540, 32'h41eaa78a} /* (10, 27, 17) {real, imag} */,
  {32'h40c392f4, 32'h00000000} /* (10, 27, 16) {real, imag} */,
  {32'hc2250540, 32'hc1eaa78a} /* (10, 27, 15) {real, imag} */,
  {32'h40c646e0, 32'h4298eb06} /* (10, 27, 14) {real, imag} */,
  {32'h426f91b5, 32'h42edab30} /* (10, 27, 13) {real, imag} */,
  {32'h412e6489, 32'h4282bd20} /* (10, 27, 12) {real, imag} */,
  {32'h42a2a73e, 32'hc2eed5b0} /* (10, 27, 11) {real, imag} */,
  {32'h41c44317, 32'hc23ab8b9} /* (10, 27, 10) {real, imag} */,
  {32'hc29cb432, 32'hc2ebbdfe} /* (10, 27, 9) {real, imag} */,
  {32'hc155a0d0, 32'hc2825c40} /* (10, 27, 8) {real, imag} */,
  {32'h4334948d, 32'h42a244dd} /* (10, 27, 7) {real, imag} */,
  {32'h40afeb08, 32'hc181215d} /* (10, 27, 6) {real, imag} */,
  {32'hc3165064, 32'h4190605c} /* (10, 27, 5) {real, imag} */,
  {32'h42c3923a, 32'h42d8ce28} /* (10, 27, 4) {real, imag} */,
  {32'hc21e0849, 32'hc319e569} /* (10, 27, 3) {real, imag} */,
  {32'hc4ec8f80, 32'hc39e8ed7} /* (10, 27, 2) {real, imag} */,
  {32'h45aef8f8, 32'h448aca0f} /* (10, 27, 1) {real, imag} */,
  {32'h45b32c28, 32'h00000000} /* (10, 27, 0) {real, imag} */,
  {32'h45a79d8d, 32'hc42e7222} /* (10, 26, 31) {real, imag} */,
  {32'hc4ee9508, 32'h435d0ac0} /* (10, 26, 30) {real, imag} */,
  {32'hc1501076, 32'h42967686} /* (10, 26, 29) {real, imag} */,
  {32'h4363ce5d, 32'hc282ccf4} /* (10, 26, 28) {real, imag} */,
  {32'hc30b4066, 32'h43081f1f} /* (10, 26, 27) {real, imag} */,
  {32'hc330252b, 32'hc278af61} /* (10, 26, 26) {real, imag} */,
  {32'h413947d4, 32'h42375f27} /* (10, 26, 25) {real, imag} */,
  {32'hc300488f, 32'h42dc4bbf} /* (10, 26, 24) {real, imag} */,
  {32'h42dde07c, 32'h425ab044} /* (10, 26, 23) {real, imag} */,
  {32'hc20b4f65, 32'hc290e732} /* (10, 26, 22) {real, imag} */,
  {32'h4121c2cc, 32'h41aea934} /* (10, 26, 21) {real, imag} */,
  {32'h428b5b5f, 32'h41450dc0} /* (10, 26, 20) {real, imag} */,
  {32'h42d65b86, 32'hc303cc95} /* (10, 26, 19) {real, imag} */,
  {32'h4280628e, 32'hc2d2881f} /* (10, 26, 18) {real, imag} */,
  {32'hc1d67ac8, 32'h42216e96} /* (10, 26, 17) {real, imag} */,
  {32'hc28b3b5c, 32'h00000000} /* (10, 26, 16) {real, imag} */,
  {32'hc1d67ac8, 32'hc2216e96} /* (10, 26, 15) {real, imag} */,
  {32'h4280628e, 32'h42d2881f} /* (10, 26, 14) {real, imag} */,
  {32'h42d65b86, 32'h4303cc95} /* (10, 26, 13) {real, imag} */,
  {32'h428b5b5f, 32'hc1450dc0} /* (10, 26, 12) {real, imag} */,
  {32'h4121c2cc, 32'hc1aea934} /* (10, 26, 11) {real, imag} */,
  {32'hc20b4f65, 32'h4290e732} /* (10, 26, 10) {real, imag} */,
  {32'h42dde07c, 32'hc25ab044} /* (10, 26, 9) {real, imag} */,
  {32'hc300488f, 32'hc2dc4bbf} /* (10, 26, 8) {real, imag} */,
  {32'h413947d4, 32'hc2375f27} /* (10, 26, 7) {real, imag} */,
  {32'hc330252b, 32'h4278af61} /* (10, 26, 6) {real, imag} */,
  {32'hc30b4066, 32'hc3081f1f} /* (10, 26, 5) {real, imag} */,
  {32'h4363ce5d, 32'h4282ccf4} /* (10, 26, 4) {real, imag} */,
  {32'hc1501076, 32'hc2967686} /* (10, 26, 3) {real, imag} */,
  {32'hc4ee9508, 32'hc35d0ac0} /* (10, 26, 2) {real, imag} */,
  {32'h45a79d8d, 32'h442e7222} /* (10, 26, 1) {real, imag} */,
  {32'h45a8b93b, 32'h00000000} /* (10, 26, 0) {real, imag} */,
  {32'h4599a6c9, 32'hc3c91c94} /* (10, 25, 31) {real, imag} */,
  {32'hc4e887b2, 32'h4396e2dc} /* (10, 25, 30) {real, imag} */,
  {32'hc2129858, 32'h4184f95e} /* (10, 25, 29) {real, imag} */,
  {32'h42eb3ff6, 32'hc2e1978c} /* (10, 25, 28) {real, imag} */,
  {32'hc2be79c8, 32'h42a45232} /* (10, 25, 27) {real, imag} */,
  {32'hc26c63bd, 32'hc2b1df4d} /* (10, 25, 26) {real, imag} */,
  {32'h403b9738, 32'h428f136e} /* (10, 25, 25) {real, imag} */,
  {32'h4190ffd9, 32'h42cbde30} /* (10, 25, 24) {real, imag} */,
  {32'h42924226, 32'h42415bef} /* (10, 25, 23) {real, imag} */,
  {32'hc1ca6bac, 32'hc2ca50ec} /* (10, 25, 22) {real, imag} */,
  {32'hc264e0aa, 32'hc1a03d7f} /* (10, 25, 21) {real, imag} */,
  {32'hc2246f26, 32'hc22fa6b8} /* (10, 25, 20) {real, imag} */,
  {32'hc1500a6d, 32'h423811b4} /* (10, 25, 19) {real, imag} */,
  {32'hc1dcae1c, 32'hc2999d88} /* (10, 25, 18) {real, imag} */,
  {32'hc24498c7, 32'h413add78} /* (10, 25, 17) {real, imag} */,
  {32'hc15710a8, 32'h00000000} /* (10, 25, 16) {real, imag} */,
  {32'hc24498c7, 32'hc13add78} /* (10, 25, 15) {real, imag} */,
  {32'hc1dcae1c, 32'h42999d88} /* (10, 25, 14) {real, imag} */,
  {32'hc1500a6d, 32'hc23811b4} /* (10, 25, 13) {real, imag} */,
  {32'hc2246f26, 32'h422fa6b8} /* (10, 25, 12) {real, imag} */,
  {32'hc264e0aa, 32'h41a03d7f} /* (10, 25, 11) {real, imag} */,
  {32'hc1ca6bac, 32'h42ca50ec} /* (10, 25, 10) {real, imag} */,
  {32'h42924226, 32'hc2415bef} /* (10, 25, 9) {real, imag} */,
  {32'h4190ffd9, 32'hc2cbde30} /* (10, 25, 8) {real, imag} */,
  {32'h403b9738, 32'hc28f136e} /* (10, 25, 7) {real, imag} */,
  {32'hc26c63bd, 32'h42b1df4d} /* (10, 25, 6) {real, imag} */,
  {32'hc2be79c8, 32'hc2a45232} /* (10, 25, 5) {real, imag} */,
  {32'h42eb3ff6, 32'h42e1978c} /* (10, 25, 4) {real, imag} */,
  {32'hc2129858, 32'hc184f95e} /* (10, 25, 3) {real, imag} */,
  {32'hc4e887b2, 32'hc396e2dc} /* (10, 25, 2) {real, imag} */,
  {32'h4599a6c9, 32'h43c91c94} /* (10, 25, 1) {real, imag} */,
  {32'h45994bc2, 32'h00000000} /* (10, 25, 0) {real, imag} */,
  {32'h45895a36, 32'hc36b3350} /* (10, 24, 31) {real, imag} */,
  {32'hc4c23e0f, 32'h434da510} /* (10, 24, 30) {real, imag} */,
  {32'hc3408e56, 32'h3ebcdf80} /* (10, 24, 29) {real, imag} */,
  {32'h4381845a, 32'hc1e7a988} /* (10, 24, 28) {real, imag} */,
  {32'hc33d0116, 32'h43694a81} /* (10, 24, 27) {real, imag} */,
  {32'hc2a90ecc, 32'h42adb81a} /* (10, 24, 26) {real, imag} */,
  {32'h428c68a6, 32'hbff9d600} /* (10, 24, 25) {real, imag} */,
  {32'hc2f28647, 32'h42260cfa} /* (10, 24, 24) {real, imag} */,
  {32'h424072b3, 32'hc2678f7a} /* (10, 24, 23) {real, imag} */,
  {32'h4281791a, 32'hc2806e7d} /* (10, 24, 22) {real, imag} */,
  {32'hc2955b6d, 32'h425dcbff} /* (10, 24, 21) {real, imag} */,
  {32'h4291c43f, 32'hc2c4efb3} /* (10, 24, 20) {real, imag} */,
  {32'h4251654a, 32'hc1ab9638} /* (10, 24, 19) {real, imag} */,
  {32'h4298a3f8, 32'hc116e584} /* (10, 24, 18) {real, imag} */,
  {32'h429f6c5e, 32'hc28790a5} /* (10, 24, 17) {real, imag} */,
  {32'h4240a552, 32'h00000000} /* (10, 24, 16) {real, imag} */,
  {32'h429f6c5e, 32'h428790a5} /* (10, 24, 15) {real, imag} */,
  {32'h4298a3f8, 32'h4116e584} /* (10, 24, 14) {real, imag} */,
  {32'h4251654a, 32'h41ab9638} /* (10, 24, 13) {real, imag} */,
  {32'h4291c43f, 32'h42c4efb3} /* (10, 24, 12) {real, imag} */,
  {32'hc2955b6d, 32'hc25dcbff} /* (10, 24, 11) {real, imag} */,
  {32'h4281791a, 32'h42806e7d} /* (10, 24, 10) {real, imag} */,
  {32'h424072b3, 32'h42678f7a} /* (10, 24, 9) {real, imag} */,
  {32'hc2f28647, 32'hc2260cfa} /* (10, 24, 8) {real, imag} */,
  {32'h428c68a6, 32'h3ff9d600} /* (10, 24, 7) {real, imag} */,
  {32'hc2a90ecc, 32'hc2adb81a} /* (10, 24, 6) {real, imag} */,
  {32'hc33d0116, 32'hc3694a81} /* (10, 24, 5) {real, imag} */,
  {32'h4381845a, 32'h41e7a988} /* (10, 24, 4) {real, imag} */,
  {32'hc3408e56, 32'hbebcdf80} /* (10, 24, 3) {real, imag} */,
  {32'hc4c23e0f, 32'hc34da510} /* (10, 24, 2) {real, imag} */,
  {32'h45895a36, 32'h436b3350} /* (10, 24, 1) {real, imag} */,
  {32'h45851561, 32'h00000000} /* (10, 24, 0) {real, imag} */,
  {32'h455dafa0, 32'hc2101ee0} /* (10, 23, 31) {real, imag} */,
  {32'hc4a45294, 32'h43055d0a} /* (10, 23, 30) {real, imag} */,
  {32'hc3643eb2, 32'h42f1491d} /* (10, 23, 29) {real, imag} */,
  {32'h43a2a212, 32'hc30fccd7} /* (10, 23, 28) {real, imag} */,
  {32'hc35bb39b, 32'h439c1384} /* (10, 23, 27) {real, imag} */,
  {32'hc17a2eec, 32'hc1c89022} /* (10, 23, 26) {real, imag} */,
  {32'h40e1f5d0, 32'hc0526a60} /* (10, 23, 25) {real, imag} */,
  {32'hc2a9c799, 32'h43092064} /* (10, 23, 24) {real, imag} */,
  {32'h428b313e, 32'hc2168ac4} /* (10, 23, 23) {real, imag} */,
  {32'h42b271db, 32'hc29a0eca} /* (10, 23, 22) {real, imag} */,
  {32'hc194509d, 32'h431f4596} /* (10, 23, 21) {real, imag} */,
  {32'h42317465, 32'h42640eb8} /* (10, 23, 20) {real, imag} */,
  {32'hc298e2bf, 32'hc28ac306} /* (10, 23, 19) {real, imag} */,
  {32'hc206dc6f, 32'h4213096f} /* (10, 23, 18) {real, imag} */,
  {32'hc0241628, 32'h4187fd3c} /* (10, 23, 17) {real, imag} */,
  {32'hbd0e3400, 32'h00000000} /* (10, 23, 16) {real, imag} */,
  {32'hc0241628, 32'hc187fd3c} /* (10, 23, 15) {real, imag} */,
  {32'hc206dc6f, 32'hc213096f} /* (10, 23, 14) {real, imag} */,
  {32'hc298e2bf, 32'h428ac306} /* (10, 23, 13) {real, imag} */,
  {32'h42317465, 32'hc2640eb8} /* (10, 23, 12) {real, imag} */,
  {32'hc194509d, 32'hc31f4596} /* (10, 23, 11) {real, imag} */,
  {32'h42b271db, 32'h429a0eca} /* (10, 23, 10) {real, imag} */,
  {32'h428b313e, 32'h42168ac4} /* (10, 23, 9) {real, imag} */,
  {32'hc2a9c799, 32'hc3092064} /* (10, 23, 8) {real, imag} */,
  {32'h40e1f5d0, 32'h40526a60} /* (10, 23, 7) {real, imag} */,
  {32'hc17a2eec, 32'h41c89022} /* (10, 23, 6) {real, imag} */,
  {32'hc35bb39b, 32'hc39c1384} /* (10, 23, 5) {real, imag} */,
  {32'h43a2a212, 32'h430fccd7} /* (10, 23, 4) {real, imag} */,
  {32'hc3643eb2, 32'hc2f1491d} /* (10, 23, 3) {real, imag} */,
  {32'hc4a45294, 32'hc3055d0a} /* (10, 23, 2) {real, imag} */,
  {32'h455dafa0, 32'h42101ee0} /* (10, 23, 1) {real, imag} */,
  {32'h45513cf4, 32'h00000000} /* (10, 23, 0) {real, imag} */,
  {32'h451b0e92, 32'hc2e9904c} /* (10, 22, 31) {real, imag} */,
  {32'hc45220f2, 32'h42ec1e2a} /* (10, 22, 30) {real, imag} */,
  {32'hc30230c2, 32'h43156bd6} /* (10, 22, 29) {real, imag} */,
  {32'h433bbb67, 32'hc1a4e6dc} /* (10, 22, 28) {real, imag} */,
  {32'hc351dee8, 32'h428a42ca} /* (10, 22, 27) {real, imag} */,
  {32'h42c44452, 32'h4265f7f0} /* (10, 22, 26) {real, imag} */,
  {32'hc3361fde, 32'hc1bfdf74} /* (10, 22, 25) {real, imag} */,
  {32'hc28c0b40, 32'h4251a38e} /* (10, 22, 24) {real, imag} */,
  {32'hc0aca9dc, 32'hbf950aa0} /* (10, 22, 23) {real, imag} */,
  {32'hc2015257, 32'hc2dd64e8} /* (10, 22, 22) {real, imag} */,
  {32'h41c22396, 32'h41745ec9} /* (10, 22, 21) {real, imag} */,
  {32'hc263b494, 32'hc274ca72} /* (10, 22, 20) {real, imag} */,
  {32'h4208746d, 32'h4143b09c} /* (10, 22, 19) {real, imag} */,
  {32'h42677ef1, 32'h428a8378} /* (10, 22, 18) {real, imag} */,
  {32'h422d3d70, 32'hc095ad94} /* (10, 22, 17) {real, imag} */,
  {32'h42af7758, 32'h00000000} /* (10, 22, 16) {real, imag} */,
  {32'h422d3d70, 32'h4095ad94} /* (10, 22, 15) {real, imag} */,
  {32'h42677ef1, 32'hc28a8378} /* (10, 22, 14) {real, imag} */,
  {32'h4208746d, 32'hc143b09c} /* (10, 22, 13) {real, imag} */,
  {32'hc263b494, 32'h4274ca72} /* (10, 22, 12) {real, imag} */,
  {32'h41c22396, 32'hc1745ec9} /* (10, 22, 11) {real, imag} */,
  {32'hc2015257, 32'h42dd64e8} /* (10, 22, 10) {real, imag} */,
  {32'hc0aca9dc, 32'h3f950aa0} /* (10, 22, 9) {real, imag} */,
  {32'hc28c0b40, 32'hc251a38e} /* (10, 22, 8) {real, imag} */,
  {32'hc3361fde, 32'h41bfdf74} /* (10, 22, 7) {real, imag} */,
  {32'h42c44452, 32'hc265f7f0} /* (10, 22, 6) {real, imag} */,
  {32'hc351dee8, 32'hc28a42ca} /* (10, 22, 5) {real, imag} */,
  {32'h433bbb67, 32'h41a4e6dc} /* (10, 22, 4) {real, imag} */,
  {32'hc30230c2, 32'hc3156bd6} /* (10, 22, 3) {real, imag} */,
  {32'hc45220f2, 32'hc2ec1e2a} /* (10, 22, 2) {real, imag} */,
  {32'h451b0e92, 32'h42e9904c} /* (10, 22, 1) {real, imag} */,
  {32'h450afd88, 32'h00000000} /* (10, 22, 0) {real, imag} */,
  {32'h442f3040, 32'hc2b83a24} /* (10, 21, 31) {real, imag} */,
  {32'hc33bd36e, 32'hc03b7980} /* (10, 21, 30) {real, imag} */,
  {32'hc1c4880e, 32'h4298e9de} /* (10, 21, 29) {real, imag} */,
  {32'h42b75536, 32'hc28a7289} /* (10, 21, 28) {real, imag} */,
  {32'hc33c9fc6, 32'h421fadc2} /* (10, 21, 27) {real, imag} */,
  {32'h42e8524c, 32'h41930bf7} /* (10, 21, 26) {real, imag} */,
  {32'hc1e72246, 32'hc28c6292} /* (10, 21, 25) {real, imag} */,
  {32'hc2836b6a, 32'h42615fc0} /* (10, 21, 24) {real, imag} */,
  {32'hc25a140c, 32'h4291def4} /* (10, 21, 23) {real, imag} */,
  {32'hc23049aa, 32'hc20585cf} /* (10, 21, 22) {real, imag} */,
  {32'h42151d41, 32'h42a6bc14} /* (10, 21, 21) {real, imag} */,
  {32'h429b72e7, 32'hc22ff6dd} /* (10, 21, 20) {real, imag} */,
  {32'h421735af, 32'h422d2411} /* (10, 21, 19) {real, imag} */,
  {32'h423b73ee, 32'hc0f01afa} /* (10, 21, 18) {real, imag} */,
  {32'h426da5be, 32'h41d4e52e} /* (10, 21, 17) {real, imag} */,
  {32'hc129c02a, 32'h00000000} /* (10, 21, 16) {real, imag} */,
  {32'h426da5be, 32'hc1d4e52e} /* (10, 21, 15) {real, imag} */,
  {32'h423b73ee, 32'h40f01afa} /* (10, 21, 14) {real, imag} */,
  {32'h421735af, 32'hc22d2411} /* (10, 21, 13) {real, imag} */,
  {32'h429b72e7, 32'h422ff6dd} /* (10, 21, 12) {real, imag} */,
  {32'h42151d41, 32'hc2a6bc14} /* (10, 21, 11) {real, imag} */,
  {32'hc23049aa, 32'h420585cf} /* (10, 21, 10) {real, imag} */,
  {32'hc25a140c, 32'hc291def4} /* (10, 21, 9) {real, imag} */,
  {32'hc2836b6a, 32'hc2615fc0} /* (10, 21, 8) {real, imag} */,
  {32'hc1e72246, 32'h428c6292} /* (10, 21, 7) {real, imag} */,
  {32'h42e8524c, 32'hc1930bf7} /* (10, 21, 6) {real, imag} */,
  {32'hc33c9fc6, 32'hc21fadc2} /* (10, 21, 5) {real, imag} */,
  {32'h42b75536, 32'h428a7289} /* (10, 21, 4) {real, imag} */,
  {32'hc1c4880e, 32'hc298e9de} /* (10, 21, 3) {real, imag} */,
  {32'hc33bd36e, 32'h403b7980} /* (10, 21, 2) {real, imag} */,
  {32'h442f3040, 32'h42b83a24} /* (10, 21, 1) {real, imag} */,
  {32'h446f4988, 32'h00000000} /* (10, 21, 0) {real, imag} */,
  {32'hc4a872a6, 32'h42e724b8} /* (10, 20, 31) {real, imag} */,
  {32'h441e1a40, 32'hc3924854} /* (10, 20, 30) {real, imag} */,
  {32'hc28f0d60, 32'h40f924c0} /* (10, 20, 29) {real, imag} */,
  {32'hc34558de, 32'hc204a954} /* (10, 20, 28) {real, imag} */,
  {32'h4278acc8, 32'h42a43bbf} /* (10, 20, 27) {real, imag} */,
  {32'h42694556, 32'hc30b6ff9} /* (10, 20, 26) {real, imag} */,
  {32'h408b8f48, 32'h420e41b6} /* (10, 20, 25) {real, imag} */,
  {32'h42546e18, 32'hc20947df} /* (10, 20, 24) {real, imag} */,
  {32'hc299c178, 32'h41888b51} /* (10, 20, 23) {real, imag} */,
  {32'h41a61f23, 32'hc2101020} /* (10, 20, 22) {real, imag} */,
  {32'hc16034fa, 32'hc21cef4e} /* (10, 20, 21) {real, imag} */,
  {32'hc0a90a48, 32'hc1719544} /* (10, 20, 20) {real, imag} */,
  {32'hc2d5566c, 32'hc2b24178} /* (10, 20, 19) {real, imag} */,
  {32'h4221e2b0, 32'hc2ab0552} /* (10, 20, 18) {real, imag} */,
  {32'h42367b08, 32'hc1b7d40f} /* (10, 20, 17) {real, imag} */,
  {32'hc16c4d3e, 32'h00000000} /* (10, 20, 16) {real, imag} */,
  {32'h42367b08, 32'h41b7d40f} /* (10, 20, 15) {real, imag} */,
  {32'h4221e2b0, 32'h42ab0552} /* (10, 20, 14) {real, imag} */,
  {32'hc2d5566c, 32'h42b24178} /* (10, 20, 13) {real, imag} */,
  {32'hc0a90a48, 32'h41719544} /* (10, 20, 12) {real, imag} */,
  {32'hc16034fa, 32'h421cef4e} /* (10, 20, 11) {real, imag} */,
  {32'h41a61f23, 32'h42101020} /* (10, 20, 10) {real, imag} */,
  {32'hc299c178, 32'hc1888b51} /* (10, 20, 9) {real, imag} */,
  {32'h42546e18, 32'h420947df} /* (10, 20, 8) {real, imag} */,
  {32'h408b8f48, 32'hc20e41b6} /* (10, 20, 7) {real, imag} */,
  {32'h42694556, 32'h430b6ff9} /* (10, 20, 6) {real, imag} */,
  {32'h4278acc8, 32'hc2a43bbf} /* (10, 20, 5) {real, imag} */,
  {32'hc34558de, 32'h4204a954} /* (10, 20, 4) {real, imag} */,
  {32'hc28f0d60, 32'hc0f924c0} /* (10, 20, 3) {real, imag} */,
  {32'h441e1a40, 32'h43924854} /* (10, 20, 2) {real, imag} */,
  {32'hc4a872a6, 32'hc2e724b8} /* (10, 20, 1) {real, imag} */,
  {32'hc410e206, 32'h00000000} /* (10, 20, 0) {real, imag} */,
  {32'hc52b8027, 32'h43be2790} /* (10, 19, 31) {real, imag} */,
  {32'h4480ce54, 32'hc3ab1fcd} /* (10, 19, 30) {real, imag} */,
  {32'hc30b7e36, 32'h42a0547c} /* (10, 19, 29) {real, imag} */,
  {32'hc2abc276, 32'h42c1e131} /* (10, 19, 28) {real, imag} */,
  {32'h42e3f0d0, 32'h41b1e204} /* (10, 19, 27) {real, imag} */,
  {32'h4221af82, 32'hc27c98fa} /* (10, 19, 26) {real, imag} */,
  {32'hc2570d99, 32'h40aa0f50} /* (10, 19, 25) {real, imag} */,
  {32'h428d2829, 32'hc27e8e72} /* (10, 19, 24) {real, imag} */,
  {32'hc118e873, 32'hc2a89234} /* (10, 19, 23) {real, imag} */,
  {32'h421b403e, 32'hc1dca57c} /* (10, 19, 22) {real, imag} */,
  {32'h42945c52, 32'hc18aa892} /* (10, 19, 21) {real, imag} */,
  {32'h41956078, 32'h4210ed90} /* (10, 19, 20) {real, imag} */,
  {32'hc1e31c94, 32'h3f7195a0} /* (10, 19, 19) {real, imag} */,
  {32'hc15f1693, 32'h427de251} /* (10, 19, 18) {real, imag} */,
  {32'hc20d2002, 32'hc2889e5c} /* (10, 19, 17) {real, imag} */,
  {32'hbead69c0, 32'h00000000} /* (10, 19, 16) {real, imag} */,
  {32'hc20d2002, 32'h42889e5c} /* (10, 19, 15) {real, imag} */,
  {32'hc15f1693, 32'hc27de251} /* (10, 19, 14) {real, imag} */,
  {32'hc1e31c94, 32'hbf7195a0} /* (10, 19, 13) {real, imag} */,
  {32'h41956078, 32'hc210ed90} /* (10, 19, 12) {real, imag} */,
  {32'h42945c52, 32'h418aa892} /* (10, 19, 11) {real, imag} */,
  {32'h421b403e, 32'h41dca57c} /* (10, 19, 10) {real, imag} */,
  {32'hc118e873, 32'h42a89234} /* (10, 19, 9) {real, imag} */,
  {32'h428d2829, 32'h427e8e72} /* (10, 19, 8) {real, imag} */,
  {32'hc2570d99, 32'hc0aa0f50} /* (10, 19, 7) {real, imag} */,
  {32'h4221af82, 32'h427c98fa} /* (10, 19, 6) {real, imag} */,
  {32'h42e3f0d0, 32'hc1b1e204} /* (10, 19, 5) {real, imag} */,
  {32'hc2abc276, 32'hc2c1e131} /* (10, 19, 4) {real, imag} */,
  {32'hc30b7e36, 32'hc2a0547c} /* (10, 19, 3) {real, imag} */,
  {32'h4480ce54, 32'h43ab1fcd} /* (10, 19, 2) {real, imag} */,
  {32'hc52b8027, 32'hc3be2790} /* (10, 19, 1) {real, imag} */,
  {32'hc4e9e0f7, 32'h00000000} /* (10, 19, 0) {real, imag} */,
  {32'hc567cf78, 32'h43a3eca6} /* (10, 18, 31) {real, imag} */,
  {32'h44affd84, 32'hc3d3d923} /* (10, 18, 30) {real, imag} */,
  {32'h42ab600f, 32'h435c23f8} /* (10, 18, 29) {real, imag} */,
  {32'hc31e1ab6, 32'h4235363c} /* (10, 18, 28) {real, imag} */,
  {32'h430a0924, 32'hc2a9e1da} /* (10, 18, 27) {real, imag} */,
  {32'h42c90e8e, 32'hc231d8fe} /* (10, 18, 26) {real, imag} */,
  {32'hc28385fc, 32'h4242131a} /* (10, 18, 25) {real, imag} */,
  {32'h420a51cc, 32'h40ef9440} /* (10, 18, 24) {real, imag} */,
  {32'hc2876c10, 32'h42da33f0} /* (10, 18, 23) {real, imag} */,
  {32'h42844687, 32'hc2965f77} /* (10, 18, 22) {real, imag} */,
  {32'h430037e0, 32'hc28ebfdf} /* (10, 18, 21) {real, imag} */,
  {32'hc2850334, 32'hc1ef88b5} /* (10, 18, 20) {real, imag} */,
  {32'hc1c7499c, 32'hc242b1a6} /* (10, 18, 19) {real, imag} */,
  {32'hc13808d8, 32'hc317a3a6} /* (10, 18, 18) {real, imag} */,
  {32'hc2009f84, 32'hc216b921} /* (10, 18, 17) {real, imag} */,
  {32'hc2c4f10e, 32'h00000000} /* (10, 18, 16) {real, imag} */,
  {32'hc2009f84, 32'h4216b921} /* (10, 18, 15) {real, imag} */,
  {32'hc13808d8, 32'h4317a3a6} /* (10, 18, 14) {real, imag} */,
  {32'hc1c7499c, 32'h4242b1a6} /* (10, 18, 13) {real, imag} */,
  {32'hc2850334, 32'h41ef88b5} /* (10, 18, 12) {real, imag} */,
  {32'h430037e0, 32'h428ebfdf} /* (10, 18, 11) {real, imag} */,
  {32'h42844687, 32'h42965f77} /* (10, 18, 10) {real, imag} */,
  {32'hc2876c10, 32'hc2da33f0} /* (10, 18, 9) {real, imag} */,
  {32'h420a51cc, 32'hc0ef9440} /* (10, 18, 8) {real, imag} */,
  {32'hc28385fc, 32'hc242131a} /* (10, 18, 7) {real, imag} */,
  {32'h42c90e8e, 32'h4231d8fe} /* (10, 18, 6) {real, imag} */,
  {32'h430a0924, 32'h42a9e1da} /* (10, 18, 5) {real, imag} */,
  {32'hc31e1ab6, 32'hc235363c} /* (10, 18, 4) {real, imag} */,
  {32'h42ab600f, 32'hc35c23f8} /* (10, 18, 3) {real, imag} */,
  {32'h44affd84, 32'h43d3d923} /* (10, 18, 2) {real, imag} */,
  {32'hc567cf78, 32'hc3a3eca6} /* (10, 18, 1) {real, imag} */,
  {32'hc5324c5a, 32'h00000000} /* (10, 18, 0) {real, imag} */,
  {32'hc585e513, 32'h43b310d8} /* (10, 17, 31) {real, imag} */,
  {32'h44d83e41, 32'hc3c57f21} /* (10, 17, 30) {real, imag} */,
  {32'h4129c31c, 32'h425887cb} /* (10, 17, 29) {real, imag} */,
  {32'hc35d90ec, 32'h40008ba0} /* (10, 17, 28) {real, imag} */,
  {32'h4374a34a, 32'hc35b98f5} /* (10, 17, 27) {real, imag} */,
  {32'hc2345198, 32'hc1848e70} /* (10, 17, 26) {real, imag} */,
  {32'h42535d40, 32'hc212243e} /* (10, 17, 25) {real, imag} */,
  {32'h42cc9a53, 32'hc2a051be} /* (10, 17, 24) {real, imag} */,
  {32'h420627c6, 32'h42f22bef} /* (10, 17, 23) {real, imag} */,
  {32'hc2afe2dd, 32'h424db0b9} /* (10, 17, 22) {real, imag} */,
  {32'h4224ac32, 32'hc2930a32} /* (10, 17, 21) {real, imag} */,
  {32'hc2c26d6a, 32'h3e8e1600} /* (10, 17, 20) {real, imag} */,
  {32'hc197c075, 32'h41fed3e0} /* (10, 17, 19) {real, imag} */,
  {32'h4288a794, 32'h40a254dc} /* (10, 17, 18) {real, imag} */,
  {32'hc23dde0a, 32'h42747035} /* (10, 17, 17) {real, imag} */,
  {32'hc1d127c7, 32'h00000000} /* (10, 17, 16) {real, imag} */,
  {32'hc23dde0a, 32'hc2747035} /* (10, 17, 15) {real, imag} */,
  {32'h4288a794, 32'hc0a254dc} /* (10, 17, 14) {real, imag} */,
  {32'hc197c075, 32'hc1fed3e0} /* (10, 17, 13) {real, imag} */,
  {32'hc2c26d6a, 32'hbe8e1600} /* (10, 17, 12) {real, imag} */,
  {32'h4224ac32, 32'h42930a32} /* (10, 17, 11) {real, imag} */,
  {32'hc2afe2dd, 32'hc24db0b9} /* (10, 17, 10) {real, imag} */,
  {32'h420627c6, 32'hc2f22bef} /* (10, 17, 9) {real, imag} */,
  {32'h42cc9a53, 32'h42a051be} /* (10, 17, 8) {real, imag} */,
  {32'h42535d40, 32'h4212243e} /* (10, 17, 7) {real, imag} */,
  {32'hc2345198, 32'h41848e70} /* (10, 17, 6) {real, imag} */,
  {32'h4374a34a, 32'h435b98f5} /* (10, 17, 5) {real, imag} */,
  {32'hc35d90ec, 32'hc0008ba0} /* (10, 17, 4) {real, imag} */,
  {32'h4129c31c, 32'hc25887cb} /* (10, 17, 3) {real, imag} */,
  {32'h44d83e41, 32'h43c57f21} /* (10, 17, 2) {real, imag} */,
  {32'hc585e513, 32'hc3b310d8} /* (10, 17, 1) {real, imag} */,
  {32'hc5569797, 32'h00000000} /* (10, 17, 0) {real, imag} */,
  {32'hc58e7ff8, 32'h43c4e814} /* (10, 16, 31) {real, imag} */,
  {32'h44d476f2, 32'hc33b7824} /* (10, 16, 30) {real, imag} */,
  {32'hc1382708, 32'h418c3b1a} /* (10, 16, 29) {real, imag} */,
  {32'hc34652b7, 32'hc29149f0} /* (10, 16, 28) {real, imag} */,
  {32'h438e2f00, 32'hc32e465b} /* (10, 16, 27) {real, imag} */,
  {32'h418355ec, 32'hc29ab080} /* (10, 16, 26) {real, imag} */,
  {32'h41d7a34c, 32'hc2117aa3} /* (10, 16, 25) {real, imag} */,
  {32'h429bbe3c, 32'h41fa03fa} /* (10, 16, 24) {real, imag} */,
  {32'h42a37cd0, 32'h4159fdc6} /* (10, 16, 23) {real, imag} */,
  {32'h424c177b, 32'h41b04017} /* (10, 16, 22) {real, imag} */,
  {32'hc19a9b20, 32'hc23e82d9} /* (10, 16, 21) {real, imag} */,
  {32'h42a261e1, 32'hc1a60eb6} /* (10, 16, 20) {real, imag} */,
  {32'hc2cba40f, 32'h4120a0f1} /* (10, 16, 19) {real, imag} */,
  {32'h41b635c0, 32'h4238d194} /* (10, 16, 18) {real, imag} */,
  {32'hc160937b, 32'h42829e9c} /* (10, 16, 17) {real, imag} */,
  {32'hc2612b11, 32'h00000000} /* (10, 16, 16) {real, imag} */,
  {32'hc160937b, 32'hc2829e9c} /* (10, 16, 15) {real, imag} */,
  {32'h41b635c0, 32'hc238d194} /* (10, 16, 14) {real, imag} */,
  {32'hc2cba40f, 32'hc120a0f1} /* (10, 16, 13) {real, imag} */,
  {32'h42a261e1, 32'h41a60eb6} /* (10, 16, 12) {real, imag} */,
  {32'hc19a9b20, 32'h423e82d9} /* (10, 16, 11) {real, imag} */,
  {32'h424c177b, 32'hc1b04017} /* (10, 16, 10) {real, imag} */,
  {32'h42a37cd0, 32'hc159fdc6} /* (10, 16, 9) {real, imag} */,
  {32'h429bbe3c, 32'hc1fa03fa} /* (10, 16, 8) {real, imag} */,
  {32'h41d7a34c, 32'h42117aa3} /* (10, 16, 7) {real, imag} */,
  {32'h418355ec, 32'h429ab080} /* (10, 16, 6) {real, imag} */,
  {32'h438e2f00, 32'h432e465b} /* (10, 16, 5) {real, imag} */,
  {32'hc34652b7, 32'h429149f0} /* (10, 16, 4) {real, imag} */,
  {32'hc1382708, 32'hc18c3b1a} /* (10, 16, 3) {real, imag} */,
  {32'h44d476f2, 32'h433b7824} /* (10, 16, 2) {real, imag} */,
  {32'hc58e7ff8, 32'hc3c4e814} /* (10, 16, 1) {real, imag} */,
  {32'hc55776ad, 32'h00000000} /* (10, 16, 0) {real, imag} */,
  {32'hc58faf05, 32'h435c04a0} /* (10, 15, 31) {real, imag} */,
  {32'h44c84831, 32'hc3246806} /* (10, 15, 30) {real, imag} */,
  {32'h426a336b, 32'h40110b90} /* (10, 15, 29) {real, imag} */,
  {32'hc398a5fe, 32'hc21654f6} /* (10, 15, 28) {real, imag} */,
  {32'h4358a0da, 32'hc2fc59de} /* (10, 15, 27) {real, imag} */,
  {32'h4316f426, 32'hbf359c00} /* (10, 15, 26) {real, imag} */,
  {32'hc25d965e, 32'h419207c0} /* (10, 15, 25) {real, imag} */,
  {32'h4221b5d2, 32'h41dde882} /* (10, 15, 24) {real, imag} */,
  {32'h422cc6f2, 32'hc2b5202b} /* (10, 15, 23) {real, imag} */,
  {32'hbc83d000, 32'hc2a39a30} /* (10, 15, 22) {real, imag} */,
  {32'h42b09791, 32'h4144b97c} /* (10, 15, 21) {real, imag} */,
  {32'h3f762bc0, 32'hc1519680} /* (10, 15, 20) {real, imag} */,
  {32'h41f07015, 32'h421b4a38} /* (10, 15, 19) {real, imag} */,
  {32'h4299020c, 32'hc1f88ccb} /* (10, 15, 18) {real, imag} */,
  {32'hc2703bcc, 32'hc12d478c} /* (10, 15, 17) {real, imag} */,
  {32'hc112a8aa, 32'h00000000} /* (10, 15, 16) {real, imag} */,
  {32'hc2703bcc, 32'h412d478c} /* (10, 15, 15) {real, imag} */,
  {32'h4299020c, 32'h41f88ccb} /* (10, 15, 14) {real, imag} */,
  {32'h41f07015, 32'hc21b4a38} /* (10, 15, 13) {real, imag} */,
  {32'h3f762bc0, 32'h41519680} /* (10, 15, 12) {real, imag} */,
  {32'h42b09791, 32'hc144b97c} /* (10, 15, 11) {real, imag} */,
  {32'hbc83d000, 32'h42a39a30} /* (10, 15, 10) {real, imag} */,
  {32'h422cc6f2, 32'h42b5202b} /* (10, 15, 9) {real, imag} */,
  {32'h4221b5d2, 32'hc1dde882} /* (10, 15, 8) {real, imag} */,
  {32'hc25d965e, 32'hc19207c0} /* (10, 15, 7) {real, imag} */,
  {32'h4316f426, 32'h3f359c00} /* (10, 15, 6) {real, imag} */,
  {32'h4358a0da, 32'h42fc59de} /* (10, 15, 5) {real, imag} */,
  {32'hc398a5fe, 32'h421654f6} /* (10, 15, 4) {real, imag} */,
  {32'h426a336b, 32'hc0110b90} /* (10, 15, 3) {real, imag} */,
  {32'h44c84831, 32'h43246806} /* (10, 15, 2) {real, imag} */,
  {32'hc58faf05, 32'hc35c04a0} /* (10, 15, 1) {real, imag} */,
  {32'hc559e171, 32'h00000000} /* (10, 15, 0) {real, imag} */,
  {32'hc5845abe, 32'h43450a04} /* (10, 14, 31) {real, imag} */,
  {32'h44b32544, 32'hc356de32} /* (10, 14, 30) {real, imag} */,
  {32'h41db16ed, 32'h41aba214} /* (10, 14, 29) {real, imag} */,
  {32'hc36b6f32, 32'h4231e854} /* (10, 14, 28) {real, imag} */,
  {32'h428dabd1, 32'hc2de5ef2} /* (10, 14, 27) {real, imag} */,
  {32'h40854518, 32'h427cfd16} /* (10, 14, 26) {real, imag} */,
  {32'hc2680894, 32'hc2330f0e} /* (10, 14, 25) {real, imag} */,
  {32'hc2ae1248, 32'hc31ddc52} /* (10, 14, 24) {real, imag} */,
  {32'hc138c4d4, 32'hc2377c71} /* (10, 14, 23) {real, imag} */,
  {32'hc210eee4, 32'h42943ca7} /* (10, 14, 22) {real, imag} */,
  {32'hc240192a, 32'hc2bb1529} /* (10, 14, 21) {real, imag} */,
  {32'h42187d55, 32'hc1c322cf} /* (10, 14, 20) {real, imag} */,
  {32'h40235774, 32'hc261fe04} /* (10, 14, 19) {real, imag} */,
  {32'hc1f302c8, 32'hc285d9d0} /* (10, 14, 18) {real, imag} */,
  {32'hc15eb6da, 32'h4103eb25} /* (10, 14, 17) {real, imag} */,
  {32'hc1862f8a, 32'h00000000} /* (10, 14, 16) {real, imag} */,
  {32'hc15eb6da, 32'hc103eb25} /* (10, 14, 15) {real, imag} */,
  {32'hc1f302c8, 32'h4285d9d0} /* (10, 14, 14) {real, imag} */,
  {32'h40235774, 32'h4261fe04} /* (10, 14, 13) {real, imag} */,
  {32'h42187d55, 32'h41c322cf} /* (10, 14, 12) {real, imag} */,
  {32'hc240192a, 32'h42bb1529} /* (10, 14, 11) {real, imag} */,
  {32'hc210eee4, 32'hc2943ca7} /* (10, 14, 10) {real, imag} */,
  {32'hc138c4d4, 32'h42377c71} /* (10, 14, 9) {real, imag} */,
  {32'hc2ae1248, 32'h431ddc52} /* (10, 14, 8) {real, imag} */,
  {32'hc2680894, 32'h42330f0e} /* (10, 14, 7) {real, imag} */,
  {32'h40854518, 32'hc27cfd16} /* (10, 14, 6) {real, imag} */,
  {32'h428dabd1, 32'h42de5ef2} /* (10, 14, 5) {real, imag} */,
  {32'hc36b6f32, 32'hc231e854} /* (10, 14, 4) {real, imag} */,
  {32'h41db16ed, 32'hc1aba214} /* (10, 14, 3) {real, imag} */,
  {32'h44b32544, 32'h4356de32} /* (10, 14, 2) {real, imag} */,
  {32'hc5845abe, 32'hc3450a04} /* (10, 14, 1) {real, imag} */,
  {32'hc543bc7e, 32'h00000000} /* (10, 14, 0) {real, imag} */,
  {32'hc55f9a51, 32'h42ce24a0} /* (10, 13, 31) {real, imag} */,
  {32'h44a261c0, 32'hc34b4b2e} /* (10, 13, 30) {real, imag} */,
  {32'h42d92580, 32'hbdaf6a00} /* (10, 13, 29) {real, imag} */,
  {32'hc388563a, 32'h42d46a81} /* (10, 13, 28) {real, imag} */,
  {32'h42a33492, 32'hc31d2e9e} /* (10, 13, 27) {real, imag} */,
  {32'h4174885e, 32'hc21fac96} /* (10, 13, 26) {real, imag} */,
  {32'hc282c01c, 32'h40260d40} /* (10, 13, 25) {real, imag} */,
  {32'hc1ae7a48, 32'hc24d1e5e} /* (10, 13, 24) {real, imag} */,
  {32'hc0ab697a, 32'h421354ef} /* (10, 13, 23) {real, imag} */,
  {32'hc25f8b44, 32'hc1ef8224} /* (10, 13, 22) {real, imag} */,
  {32'hc167293c, 32'hc17fad6b} /* (10, 13, 21) {real, imag} */,
  {32'hc0bdf000, 32'hc2d08dca} /* (10, 13, 20) {real, imag} */,
  {32'hc275d7f0, 32'hc191e5dd} /* (10, 13, 19) {real, imag} */,
  {32'h41daddbe, 32'hc2161cd3} /* (10, 13, 18) {real, imag} */,
  {32'h42923537, 32'hc1f5765e} /* (10, 13, 17) {real, imag} */,
  {32'h41d293ff, 32'h00000000} /* (10, 13, 16) {real, imag} */,
  {32'h42923537, 32'h41f5765e} /* (10, 13, 15) {real, imag} */,
  {32'h41daddbe, 32'h42161cd3} /* (10, 13, 14) {real, imag} */,
  {32'hc275d7f0, 32'h4191e5dd} /* (10, 13, 13) {real, imag} */,
  {32'hc0bdf000, 32'h42d08dca} /* (10, 13, 12) {real, imag} */,
  {32'hc167293c, 32'h417fad6b} /* (10, 13, 11) {real, imag} */,
  {32'hc25f8b44, 32'h41ef8224} /* (10, 13, 10) {real, imag} */,
  {32'hc0ab697a, 32'hc21354ef} /* (10, 13, 9) {real, imag} */,
  {32'hc1ae7a48, 32'h424d1e5e} /* (10, 13, 8) {real, imag} */,
  {32'hc282c01c, 32'hc0260d40} /* (10, 13, 7) {real, imag} */,
  {32'h4174885e, 32'h421fac96} /* (10, 13, 6) {real, imag} */,
  {32'h42a33492, 32'h431d2e9e} /* (10, 13, 5) {real, imag} */,
  {32'hc388563a, 32'hc2d46a81} /* (10, 13, 4) {real, imag} */,
  {32'h42d92580, 32'h3daf6a00} /* (10, 13, 3) {real, imag} */,
  {32'h44a261c0, 32'h434b4b2e} /* (10, 13, 2) {real, imag} */,
  {32'hc55f9a51, 32'hc2ce24a0} /* (10, 13, 1) {real, imag} */,
  {32'hc51f8d68, 32'h00000000} /* (10, 13, 0) {real, imag} */,
  {32'hc5256d05, 32'hc2bfc158} /* (10, 12, 31) {real, imag} */,
  {32'h448d5cdb, 32'hc2ae932e} /* (10, 12, 30) {real, imag} */,
  {32'hc25cf89f, 32'h400ef940} /* (10, 12, 29) {real, imag} */,
  {32'hc35e849e, 32'h4331ee4f} /* (10, 12, 28) {real, imag} */,
  {32'h42da4aea, 32'h4188a16c} /* (10, 12, 27) {real, imag} */,
  {32'h41f8608d, 32'h415dfac4} /* (10, 12, 26) {real, imag} */,
  {32'hc26eeacd, 32'h40ac8754} /* (10, 12, 25) {real, imag} */,
  {32'h42ac03e2, 32'hc2096e61} /* (10, 12, 24) {real, imag} */,
  {32'hc228b8fc, 32'hc209795e} /* (10, 12, 23) {real, imag} */,
  {32'h42839d7e, 32'hc2ae3f7a} /* (10, 12, 22) {real, imag} */,
  {32'hc287331f, 32'hc2e1844d} /* (10, 12, 21) {real, imag} */,
  {32'h410520f6, 32'h42a63b44} /* (10, 12, 20) {real, imag} */,
  {32'h41adf23a, 32'hc11a4b8c} /* (10, 12, 19) {real, imag} */,
  {32'hc0d87cd0, 32'hc1fbb70a} /* (10, 12, 18) {real, imag} */,
  {32'hc106c782, 32'hc25c3f7e} /* (10, 12, 17) {real, imag} */,
  {32'hc1eedd5d, 32'h00000000} /* (10, 12, 16) {real, imag} */,
  {32'hc106c782, 32'h425c3f7e} /* (10, 12, 15) {real, imag} */,
  {32'hc0d87cd0, 32'h41fbb70a} /* (10, 12, 14) {real, imag} */,
  {32'h41adf23a, 32'h411a4b8c} /* (10, 12, 13) {real, imag} */,
  {32'h410520f6, 32'hc2a63b44} /* (10, 12, 12) {real, imag} */,
  {32'hc287331f, 32'h42e1844d} /* (10, 12, 11) {real, imag} */,
  {32'h42839d7e, 32'h42ae3f7a} /* (10, 12, 10) {real, imag} */,
  {32'hc228b8fc, 32'h4209795e} /* (10, 12, 9) {real, imag} */,
  {32'h42ac03e2, 32'h42096e61} /* (10, 12, 8) {real, imag} */,
  {32'hc26eeacd, 32'hc0ac8754} /* (10, 12, 7) {real, imag} */,
  {32'h41f8608d, 32'hc15dfac4} /* (10, 12, 6) {real, imag} */,
  {32'h42da4aea, 32'hc188a16c} /* (10, 12, 5) {real, imag} */,
  {32'hc35e849e, 32'hc331ee4f} /* (10, 12, 4) {real, imag} */,
  {32'hc25cf89f, 32'hc00ef940} /* (10, 12, 3) {real, imag} */,
  {32'h448d5cdb, 32'h42ae932e} /* (10, 12, 2) {real, imag} */,
  {32'hc5256d05, 32'h42bfc158} /* (10, 12, 1) {real, imag} */,
  {32'hc4d85a0d, 32'h00000000} /* (10, 12, 0) {real, imag} */,
  {32'hc4b4c768, 32'hc38be97f} /* (10, 11, 31) {real, imag} */,
  {32'h441ce07a, 32'hc1397220} /* (10, 11, 30) {real, imag} */,
  {32'hc265e3e9, 32'hc284fa76} /* (10, 11, 29) {real, imag} */,
  {32'hc209f2d3, 32'hc1fd806c} /* (10, 11, 28) {real, imag} */,
  {32'h4252398e, 32'hc2bc2ac7} /* (10, 11, 27) {real, imag} */,
  {32'hc20eabab, 32'hc224f818} /* (10, 11, 26) {real, imag} */,
  {32'h4123791c, 32'h425a1184} /* (10, 11, 25) {real, imag} */,
  {32'h422e737c, 32'hc2753eb6} /* (10, 11, 24) {real, imag} */,
  {32'h411ebfb0, 32'h430c30e2} /* (10, 11, 23) {real, imag} */,
  {32'hc18d1975, 32'hc118e063} /* (10, 11, 22) {real, imag} */,
  {32'h3e29b100, 32'h4202c0ed} /* (10, 11, 21) {real, imag} */,
  {32'h429445b5, 32'h41ec415a} /* (10, 11, 20) {real, imag} */,
  {32'h404acc10, 32'h41d5d1b2} /* (10, 11, 19) {real, imag} */,
  {32'h424364d8, 32'hc197fe9e} /* (10, 11, 18) {real, imag} */,
  {32'hc1bf1eb5, 32'h4257a0b7} /* (10, 11, 17) {real, imag} */,
  {32'hc2332e84, 32'h00000000} /* (10, 11, 16) {real, imag} */,
  {32'hc1bf1eb5, 32'hc257a0b7} /* (10, 11, 15) {real, imag} */,
  {32'h424364d8, 32'h4197fe9e} /* (10, 11, 14) {real, imag} */,
  {32'h404acc10, 32'hc1d5d1b2} /* (10, 11, 13) {real, imag} */,
  {32'h429445b5, 32'hc1ec415a} /* (10, 11, 12) {real, imag} */,
  {32'h3e29b100, 32'hc202c0ed} /* (10, 11, 11) {real, imag} */,
  {32'hc18d1975, 32'h4118e063} /* (10, 11, 10) {real, imag} */,
  {32'h411ebfb0, 32'hc30c30e2} /* (10, 11, 9) {real, imag} */,
  {32'h422e737c, 32'h42753eb6} /* (10, 11, 8) {real, imag} */,
  {32'h4123791c, 32'hc25a1184} /* (10, 11, 7) {real, imag} */,
  {32'hc20eabab, 32'h4224f818} /* (10, 11, 6) {real, imag} */,
  {32'h4252398e, 32'h42bc2ac7} /* (10, 11, 5) {real, imag} */,
  {32'hc209f2d3, 32'h41fd806c} /* (10, 11, 4) {real, imag} */,
  {32'hc265e3e9, 32'h4284fa76} /* (10, 11, 3) {real, imag} */,
  {32'h441ce07a, 32'h41397220} /* (10, 11, 2) {real, imag} */,
  {32'hc4b4c768, 32'h438be97f} /* (10, 11, 1) {real, imag} */,
  {32'hc322a4a0, 32'h00000000} /* (10, 11, 0) {real, imag} */,
  {32'h44061147, 32'hc424e7ae} /* (10, 10, 31) {real, imag} */,
  {32'hc39454a3, 32'h43951d3a} /* (10, 10, 30) {real, imag} */,
  {32'hc317cf4e, 32'hc2c3ab78} /* (10, 10, 29) {real, imag} */,
  {32'h3fccbd80, 32'hc383277e} /* (10, 10, 28) {real, imag} */,
  {32'hc1c828b0, 32'hc220d0bc} /* (10, 10, 27) {real, imag} */,
  {32'h41cf39c8, 32'hc122eec0} /* (10, 10, 26) {real, imag} */,
  {32'hc21416e2, 32'h416307d7} /* (10, 10, 25) {real, imag} */,
  {32'hc206d488, 32'h43066298} /* (10, 10, 24) {real, imag} */,
  {32'h427fd6d4, 32'h41df2f5a} /* (10, 10, 23) {real, imag} */,
  {32'h414ed701, 32'h431fac9c} /* (10, 10, 22) {real, imag} */,
  {32'h42bd648a, 32'h41d7fd28} /* (10, 10, 21) {real, imag} */,
  {32'hc2509e0c, 32'hc2c4da3b} /* (10, 10, 20) {real, imag} */,
  {32'hc2016c9b, 32'hc1d2531c} /* (10, 10, 19) {real, imag} */,
  {32'h415df984, 32'hc2077a34} /* (10, 10, 18) {real, imag} */,
  {32'h41c75bd9, 32'h4135b2f0} /* (10, 10, 17) {real, imag} */,
  {32'hc1e0b60a, 32'h00000000} /* (10, 10, 16) {real, imag} */,
  {32'h41c75bd9, 32'hc135b2f0} /* (10, 10, 15) {real, imag} */,
  {32'h415df984, 32'h42077a34} /* (10, 10, 14) {real, imag} */,
  {32'hc2016c9b, 32'h41d2531c} /* (10, 10, 13) {real, imag} */,
  {32'hc2509e0c, 32'h42c4da3b} /* (10, 10, 12) {real, imag} */,
  {32'h42bd648a, 32'hc1d7fd28} /* (10, 10, 11) {real, imag} */,
  {32'h414ed701, 32'hc31fac9c} /* (10, 10, 10) {real, imag} */,
  {32'h427fd6d4, 32'hc1df2f5a} /* (10, 10, 9) {real, imag} */,
  {32'hc206d488, 32'hc3066298} /* (10, 10, 8) {real, imag} */,
  {32'hc21416e2, 32'hc16307d7} /* (10, 10, 7) {real, imag} */,
  {32'h41cf39c8, 32'h4122eec0} /* (10, 10, 6) {real, imag} */,
  {32'hc1c828b0, 32'h4220d0bc} /* (10, 10, 5) {real, imag} */,
  {32'h3fccbd80, 32'h4383277e} /* (10, 10, 4) {real, imag} */,
  {32'hc317cf4e, 32'h42c3ab78} /* (10, 10, 3) {real, imag} */,
  {32'hc39454a3, 32'hc3951d3a} /* (10, 10, 2) {real, imag} */,
  {32'h44061147, 32'h4424e7ae} /* (10, 10, 1) {real, imag} */,
  {32'h44b4a774, 32'h00000000} /* (10, 10, 0) {real, imag} */,
  {32'h44fe3130, 32'hc485581f} /* (10, 9, 31) {real, imag} */,
  {32'hc462e471, 32'h43a7fb88} /* (10, 9, 30) {real, imag} */,
  {32'hc2c04645, 32'hc2793c36} /* (10, 9, 29) {real, imag} */,
  {32'hc20311b8, 32'hc3329541} /* (10, 9, 28) {real, imag} */,
  {32'hc2f62e7a, 32'h433d2cc1} /* (10, 9, 27) {real, imag} */,
  {32'hc2bbc70a, 32'h42402047} /* (10, 9, 26) {real, imag} */,
  {32'h42b196c3, 32'hc2d1e515} /* (10, 9, 25) {real, imag} */,
  {32'h42463d7a, 32'h4291b4aa} /* (10, 9, 24) {real, imag} */,
  {32'h4297365e, 32'hc328969b} /* (10, 9, 23) {real, imag} */,
  {32'h41e5c993, 32'hc169aecc} /* (10, 9, 22) {real, imag} */,
  {32'h41783d5a, 32'hc216e31a} /* (10, 9, 21) {real, imag} */,
  {32'hc2a78064, 32'h42454298} /* (10, 9, 20) {real, imag} */,
  {32'h42148a02, 32'h420df79a} /* (10, 9, 19) {real, imag} */,
  {32'hc2b2be5a, 32'h420506c9} /* (10, 9, 18) {real, imag} */,
  {32'hc227ea22, 32'h42b40e0c} /* (10, 9, 17) {real, imag} */,
  {32'hc17f2fe8, 32'h00000000} /* (10, 9, 16) {real, imag} */,
  {32'hc227ea22, 32'hc2b40e0c} /* (10, 9, 15) {real, imag} */,
  {32'hc2b2be5a, 32'hc20506c9} /* (10, 9, 14) {real, imag} */,
  {32'h42148a02, 32'hc20df79a} /* (10, 9, 13) {real, imag} */,
  {32'hc2a78064, 32'hc2454298} /* (10, 9, 12) {real, imag} */,
  {32'h41783d5a, 32'h4216e31a} /* (10, 9, 11) {real, imag} */,
  {32'h41e5c993, 32'h4169aecc} /* (10, 9, 10) {real, imag} */,
  {32'h4297365e, 32'h4328969b} /* (10, 9, 9) {real, imag} */,
  {32'h42463d7a, 32'hc291b4aa} /* (10, 9, 8) {real, imag} */,
  {32'h42b196c3, 32'h42d1e515} /* (10, 9, 7) {real, imag} */,
  {32'hc2bbc70a, 32'hc2402047} /* (10, 9, 6) {real, imag} */,
  {32'hc2f62e7a, 32'hc33d2cc1} /* (10, 9, 5) {real, imag} */,
  {32'hc20311b8, 32'h43329541} /* (10, 9, 4) {real, imag} */,
  {32'hc2c04645, 32'h42793c36} /* (10, 9, 3) {real, imag} */,
  {32'hc462e471, 32'hc3a7fb88} /* (10, 9, 2) {real, imag} */,
  {32'h44fe3130, 32'h4485581f} /* (10, 9, 1) {real, imag} */,
  {32'h4529b276, 32'h00000000} /* (10, 9, 0) {real, imag} */,
  {32'h4536dd56, 32'hc4b1cb86} /* (10, 8, 31) {real, imag} */,
  {32'hc48c4af5, 32'h4415bcd2} /* (10, 8, 30) {real, imag} */,
  {32'hc3290e9c, 32'hc2390db5} /* (10, 8, 29) {real, imag} */,
  {32'h42cc379a, 32'hc280377a} /* (10, 8, 28) {real, imag} */,
  {32'hc2bc857c, 32'h4398080c} /* (10, 8, 27) {real, imag} */,
  {32'hc2193eeb, 32'h4243c8a8} /* (10, 8, 26) {real, imag} */,
  {32'h426ac400, 32'hc235ca8c} /* (10, 8, 25) {real, imag} */,
  {32'hc11fbbb8, 32'h4234e6ea} /* (10, 8, 24) {real, imag} */,
  {32'hc2b92752, 32'h41811b65} /* (10, 8, 23) {real, imag} */,
  {32'h42ad48fc, 32'h41d59ecf} /* (10, 8, 22) {real, imag} */,
  {32'h42672e87, 32'h42e3966e} /* (10, 8, 21) {real, imag} */,
  {32'hc23dab82, 32'hbfbe80c0} /* (10, 8, 20) {real, imag} */,
  {32'h42691df2, 32'hc2c15522} /* (10, 8, 19) {real, imag} */,
  {32'h42865188, 32'hc26525cb} /* (10, 8, 18) {real, imag} */,
  {32'hc03caff0, 32'hc1ff548c} /* (10, 8, 17) {real, imag} */,
  {32'hc232ea2a, 32'h00000000} /* (10, 8, 16) {real, imag} */,
  {32'hc03caff0, 32'h41ff548c} /* (10, 8, 15) {real, imag} */,
  {32'h42865188, 32'h426525cb} /* (10, 8, 14) {real, imag} */,
  {32'h42691df2, 32'h42c15522} /* (10, 8, 13) {real, imag} */,
  {32'hc23dab82, 32'h3fbe80c0} /* (10, 8, 12) {real, imag} */,
  {32'h42672e87, 32'hc2e3966e} /* (10, 8, 11) {real, imag} */,
  {32'h42ad48fc, 32'hc1d59ecf} /* (10, 8, 10) {real, imag} */,
  {32'hc2b92752, 32'hc1811b65} /* (10, 8, 9) {real, imag} */,
  {32'hc11fbbb8, 32'hc234e6ea} /* (10, 8, 8) {real, imag} */,
  {32'h426ac400, 32'h4235ca8c} /* (10, 8, 7) {real, imag} */,
  {32'hc2193eeb, 32'hc243c8a8} /* (10, 8, 6) {real, imag} */,
  {32'hc2bc857c, 32'hc398080c} /* (10, 8, 5) {real, imag} */,
  {32'h42cc379a, 32'h4280377a} /* (10, 8, 4) {real, imag} */,
  {32'hc3290e9c, 32'h42390db5} /* (10, 8, 3) {real, imag} */,
  {32'hc48c4af5, 32'hc415bcd2} /* (10, 8, 2) {real, imag} */,
  {32'h4536dd56, 32'h44b1cb86} /* (10, 8, 1) {real, imag} */,
  {32'h45673684, 32'h00000000} /* (10, 8, 0) {real, imag} */,
  {32'h455c8472, 32'hc4ece771} /* (10, 7, 31) {real, imag} */,
  {32'hc48a94ce, 32'h4453c128} /* (10, 7, 30) {real, imag} */,
  {32'hc2ffcb12, 32'hc2a966fe} /* (10, 7, 29) {real, imag} */,
  {32'h4215c80c, 32'hc30d24b1} /* (10, 7, 28) {real, imag} */,
  {32'hc2dac2a0, 32'h43541cef} /* (10, 7, 27) {real, imag} */,
  {32'hc2ced70e, 32'h42b7423d} /* (10, 7, 26) {real, imag} */,
  {32'hc0b63acc, 32'hc2153db0} /* (10, 7, 25) {real, imag} */,
  {32'hc1dbd001, 32'hc149ed94} /* (10, 7, 24) {real, imag} */,
  {32'h4252c1ab, 32'h41a6fa82} /* (10, 7, 23) {real, imag} */,
  {32'h43085b3e, 32'h42e2db70} /* (10, 7, 22) {real, imag} */,
  {32'hc1e0fefd, 32'h424c70b2} /* (10, 7, 21) {real, imag} */,
  {32'h41c3ccbc, 32'h410227a6} /* (10, 7, 20) {real, imag} */,
  {32'h40384a1c, 32'hc235efc6} /* (10, 7, 19) {real, imag} */,
  {32'hc30c1a1c, 32'h3f96c6a0} /* (10, 7, 18) {real, imag} */,
  {32'hc2768931, 32'hc19c0be8} /* (10, 7, 17) {real, imag} */,
  {32'hc2c5834b, 32'h00000000} /* (10, 7, 16) {real, imag} */,
  {32'hc2768931, 32'h419c0be8} /* (10, 7, 15) {real, imag} */,
  {32'hc30c1a1c, 32'hbf96c6a0} /* (10, 7, 14) {real, imag} */,
  {32'h40384a1c, 32'h4235efc6} /* (10, 7, 13) {real, imag} */,
  {32'h41c3ccbc, 32'hc10227a6} /* (10, 7, 12) {real, imag} */,
  {32'hc1e0fefd, 32'hc24c70b2} /* (10, 7, 11) {real, imag} */,
  {32'h43085b3e, 32'hc2e2db70} /* (10, 7, 10) {real, imag} */,
  {32'h4252c1ab, 32'hc1a6fa82} /* (10, 7, 9) {real, imag} */,
  {32'hc1dbd001, 32'h4149ed94} /* (10, 7, 8) {real, imag} */,
  {32'hc0b63acc, 32'h42153db0} /* (10, 7, 7) {real, imag} */,
  {32'hc2ced70e, 32'hc2b7423d} /* (10, 7, 6) {real, imag} */,
  {32'hc2dac2a0, 32'hc3541cef} /* (10, 7, 5) {real, imag} */,
  {32'h4215c80c, 32'h430d24b1} /* (10, 7, 4) {real, imag} */,
  {32'hc2ffcb12, 32'h42a966fe} /* (10, 7, 3) {real, imag} */,
  {32'hc48a94ce, 32'hc453c128} /* (10, 7, 2) {real, imag} */,
  {32'h455c8472, 32'h44ece771} /* (10, 7, 1) {real, imag} */,
  {32'h458d9ada, 32'h00000000} /* (10, 7, 0) {real, imag} */,
  {32'h4567af3a, 32'hc51b0e78} /* (10, 6, 31) {real, imag} */,
  {32'hc45349f4, 32'h44813d6b} /* (10, 6, 30) {real, imag} */,
  {32'hc1dbe2e5, 32'h4212284d} /* (10, 6, 29) {real, imag} */,
  {32'hc19b5938, 32'h420cf8c4} /* (10, 6, 28) {real, imag} */,
  {32'hc2d0c6c1, 32'h42db88be} /* (10, 6, 27) {real, imag} */,
  {32'h425478e4, 32'hc09e8d98} /* (10, 6, 26) {real, imag} */,
  {32'h423d75ff, 32'hc0a67198} /* (10, 6, 25) {real, imag} */,
  {32'hc11c7490, 32'hc085c8d0} /* (10, 6, 24) {real, imag} */,
  {32'h42875360, 32'hc2ab8772} /* (10, 6, 23) {real, imag} */,
  {32'h4206aabf, 32'h3fd6f9c0} /* (10, 6, 22) {real, imag} */,
  {32'hc1bb0426, 32'h4294449c} /* (10, 6, 21) {real, imag} */,
  {32'hc09acab0, 32'hc212c77a} /* (10, 6, 20) {real, imag} */,
  {32'hc050a8f0, 32'h40ef1fa0} /* (10, 6, 19) {real, imag} */,
  {32'hc2ac0f00, 32'h428d2c27} /* (10, 6, 18) {real, imag} */,
  {32'h4192b702, 32'h416e799f} /* (10, 6, 17) {real, imag} */,
  {32'hc2699bc0, 32'h00000000} /* (10, 6, 16) {real, imag} */,
  {32'h4192b702, 32'hc16e799f} /* (10, 6, 15) {real, imag} */,
  {32'hc2ac0f00, 32'hc28d2c27} /* (10, 6, 14) {real, imag} */,
  {32'hc050a8f0, 32'hc0ef1fa0} /* (10, 6, 13) {real, imag} */,
  {32'hc09acab0, 32'h4212c77a} /* (10, 6, 12) {real, imag} */,
  {32'hc1bb0426, 32'hc294449c} /* (10, 6, 11) {real, imag} */,
  {32'h4206aabf, 32'hbfd6f9c0} /* (10, 6, 10) {real, imag} */,
  {32'h42875360, 32'h42ab8772} /* (10, 6, 9) {real, imag} */,
  {32'hc11c7490, 32'h4085c8d0} /* (10, 6, 8) {real, imag} */,
  {32'h423d75ff, 32'h40a67198} /* (10, 6, 7) {real, imag} */,
  {32'h425478e4, 32'h409e8d98} /* (10, 6, 6) {real, imag} */,
  {32'hc2d0c6c1, 32'hc2db88be} /* (10, 6, 5) {real, imag} */,
  {32'hc19b5938, 32'hc20cf8c4} /* (10, 6, 4) {real, imag} */,
  {32'hc1dbe2e5, 32'hc212284d} /* (10, 6, 3) {real, imag} */,
  {32'hc45349f4, 32'hc4813d6b} /* (10, 6, 2) {real, imag} */,
  {32'h4567af3a, 32'h451b0e78} /* (10, 6, 1) {real, imag} */,
  {32'h45a09f19, 32'h00000000} /* (10, 6, 0) {real, imag} */,
  {32'h45599ed3, 32'hc54b7a08} /* (10, 5, 31) {real, imag} */,
  {32'hc3ded632, 32'h4494388f} /* (10, 5, 30) {real, imag} */,
  {32'hc2fc3d0c, 32'hc185c088} /* (10, 5, 29) {real, imag} */,
  {32'hbfbd8aa0, 32'h435883b0} /* (10, 5, 28) {real, imag} */,
  {32'hc2f663c9, 32'h435fa416} /* (10, 5, 27) {real, imag} */,
  {32'h424ae169, 32'hc1d601c7} /* (10, 5, 26) {real, imag} */,
  {32'h41a16208, 32'hc1e17894} /* (10, 5, 25) {real, imag} */,
  {32'hc2a21ae4, 32'h43178d3a} /* (10, 5, 24) {real, imag} */,
  {32'hc2cc7c32, 32'hc1fb253a} /* (10, 5, 23) {real, imag} */,
  {32'h4181c9e9, 32'h42b23cb6} /* (10, 5, 22) {real, imag} */,
  {32'hc2bb0962, 32'hc15cfefc} /* (10, 5, 21) {real, imag} */,
  {32'hc1833020, 32'hc200c51d} /* (10, 5, 20) {real, imag} */,
  {32'h4229200f, 32'h41928c12} /* (10, 5, 19) {real, imag} */,
  {32'h4231e00e, 32'h4162b9c4} /* (10, 5, 18) {real, imag} */,
  {32'hc131e263, 32'hc2a52c1c} /* (10, 5, 17) {real, imag} */,
  {32'hc276b446, 32'h00000000} /* (10, 5, 16) {real, imag} */,
  {32'hc131e263, 32'h42a52c1c} /* (10, 5, 15) {real, imag} */,
  {32'h4231e00e, 32'hc162b9c4} /* (10, 5, 14) {real, imag} */,
  {32'h4229200f, 32'hc1928c12} /* (10, 5, 13) {real, imag} */,
  {32'hc1833020, 32'h4200c51d} /* (10, 5, 12) {real, imag} */,
  {32'hc2bb0962, 32'h415cfefc} /* (10, 5, 11) {real, imag} */,
  {32'h4181c9e9, 32'hc2b23cb6} /* (10, 5, 10) {real, imag} */,
  {32'hc2cc7c32, 32'h41fb253a} /* (10, 5, 9) {real, imag} */,
  {32'hc2a21ae4, 32'hc3178d3a} /* (10, 5, 8) {real, imag} */,
  {32'h41a16208, 32'h41e17894} /* (10, 5, 7) {real, imag} */,
  {32'h424ae169, 32'h41d601c7} /* (10, 5, 6) {real, imag} */,
  {32'hc2f663c9, 32'hc35fa416} /* (10, 5, 5) {real, imag} */,
  {32'hbfbd8aa0, 32'hc35883b0} /* (10, 5, 4) {real, imag} */,
  {32'hc2fc3d0c, 32'h4185c088} /* (10, 5, 3) {real, imag} */,
  {32'hc3ded632, 32'hc494388f} /* (10, 5, 2) {real, imag} */,
  {32'h45599ed3, 32'h454b7a08} /* (10, 5, 1) {real, imag} */,
  {32'h45adf68c, 32'h00000000} /* (10, 5, 0) {real, imag} */,
  {32'h45533099, 32'hc56a8f63} /* (10, 4, 31) {real, imag} */,
  {32'hc1004e80, 32'h44938523} /* (10, 4, 30) {real, imag} */,
  {32'hc2d5bd80, 32'h40884890} /* (10, 4, 29) {real, imag} */,
  {32'hc2a4cf24, 32'h437ab093} /* (10, 4, 28) {real, imag} */,
  {32'hc2e5032a, 32'h42c61b3d} /* (10, 4, 27) {real, imag} */,
  {32'h426a5648, 32'h4259dfd9} /* (10, 4, 26) {real, imag} */,
  {32'h424aca35, 32'hc2b64626} /* (10, 4, 25) {real, imag} */,
  {32'hc2a7c35f, 32'h434902c2} /* (10, 4, 24) {real, imag} */,
  {32'hc17cf468, 32'hc2a8346c} /* (10, 4, 23) {real, imag} */,
  {32'h3ec10420, 32'h42c715f7} /* (10, 4, 22) {real, imag} */,
  {32'hc1ea7031, 32'hc234f119} /* (10, 4, 21) {real, imag} */,
  {32'hc1869b3e, 32'h429ad18a} /* (10, 4, 20) {real, imag} */,
  {32'hbe9b9040, 32'hc20cfd50} /* (10, 4, 19) {real, imag} */,
  {32'h41e7ef98, 32'h422c3576} /* (10, 4, 18) {real, imag} */,
  {32'hc23302ae, 32'h40e504a8} /* (10, 4, 17) {real, imag} */,
  {32'h414eaec4, 32'h00000000} /* (10, 4, 16) {real, imag} */,
  {32'hc23302ae, 32'hc0e504a8} /* (10, 4, 15) {real, imag} */,
  {32'h41e7ef98, 32'hc22c3576} /* (10, 4, 14) {real, imag} */,
  {32'hbe9b9040, 32'h420cfd50} /* (10, 4, 13) {real, imag} */,
  {32'hc1869b3e, 32'hc29ad18a} /* (10, 4, 12) {real, imag} */,
  {32'hc1ea7031, 32'h4234f119} /* (10, 4, 11) {real, imag} */,
  {32'h3ec10420, 32'hc2c715f7} /* (10, 4, 10) {real, imag} */,
  {32'hc17cf468, 32'h42a8346c} /* (10, 4, 9) {real, imag} */,
  {32'hc2a7c35f, 32'hc34902c2} /* (10, 4, 8) {real, imag} */,
  {32'h424aca35, 32'h42b64626} /* (10, 4, 7) {real, imag} */,
  {32'h426a5648, 32'hc259dfd9} /* (10, 4, 6) {real, imag} */,
  {32'hc2e5032a, 32'hc2c61b3d} /* (10, 4, 5) {real, imag} */,
  {32'hc2a4cf24, 32'hc37ab093} /* (10, 4, 4) {real, imag} */,
  {32'hc2d5bd80, 32'hc0884890} /* (10, 4, 3) {real, imag} */,
  {32'hc1004e80, 32'hc4938523} /* (10, 4, 2) {real, imag} */,
  {32'h45533099, 32'h456a8f63} /* (10, 4, 1) {real, imag} */,
  {32'h45b6f506, 32'h00000000} /* (10, 4, 0) {real, imag} */,
  {32'h4552a8e4, 32'hc57ff964} /* (10, 3, 31) {real, imag} */,
  {32'h436e834c, 32'h449cea44} /* (10, 3, 30) {real, imag} */,
  {32'hc16135b0, 32'h4302421e} /* (10, 3, 29) {real, imag} */,
  {32'hc32e6d5c, 32'h4392d0dc} /* (10, 3, 28) {real, imag} */,
  {32'hc33d53f2, 32'hc2853614} /* (10, 3, 27) {real, imag} */,
  {32'hc284b8f0, 32'h4259c730} /* (10, 3, 26) {real, imag} */,
  {32'h410ff9f9, 32'h422f6c11} /* (10, 3, 25) {real, imag} */,
  {32'h42f0ffc6, 32'h4314dfe1} /* (10, 3, 24) {real, imag} */,
  {32'hc1b68718, 32'hc30773f5} /* (10, 3, 23) {real, imag} */,
  {32'hc211807f, 32'hc0c6fbe0} /* (10, 3, 22) {real, imag} */,
  {32'hc06dda58, 32'h42a95434} /* (10, 3, 21) {real, imag} */,
  {32'hc2574df8, 32'h3f401df0} /* (10, 3, 20) {real, imag} */,
  {32'hc22f3fde, 32'hc2af7991} /* (10, 3, 19) {real, imag} */,
  {32'hc17d2a86, 32'h42a1a2e0} /* (10, 3, 18) {real, imag} */,
  {32'h42b4e5bc, 32'h4166073c} /* (10, 3, 17) {real, imag} */,
  {32'h4313a2dc, 32'h00000000} /* (10, 3, 16) {real, imag} */,
  {32'h42b4e5bc, 32'hc166073c} /* (10, 3, 15) {real, imag} */,
  {32'hc17d2a86, 32'hc2a1a2e0} /* (10, 3, 14) {real, imag} */,
  {32'hc22f3fde, 32'h42af7991} /* (10, 3, 13) {real, imag} */,
  {32'hc2574df8, 32'hbf401df0} /* (10, 3, 12) {real, imag} */,
  {32'hc06dda58, 32'hc2a95434} /* (10, 3, 11) {real, imag} */,
  {32'hc211807f, 32'h40c6fbe0} /* (10, 3, 10) {real, imag} */,
  {32'hc1b68718, 32'h430773f5} /* (10, 3, 9) {real, imag} */,
  {32'h42f0ffc6, 32'hc314dfe1} /* (10, 3, 8) {real, imag} */,
  {32'h410ff9f9, 32'hc22f6c11} /* (10, 3, 7) {real, imag} */,
  {32'hc284b8f0, 32'hc259c730} /* (10, 3, 6) {real, imag} */,
  {32'hc33d53f2, 32'h42853614} /* (10, 3, 5) {real, imag} */,
  {32'hc32e6d5c, 32'hc392d0dc} /* (10, 3, 4) {real, imag} */,
  {32'hc16135b0, 32'hc302421e} /* (10, 3, 3) {real, imag} */,
  {32'h436e834c, 32'hc49cea44} /* (10, 3, 2) {real, imag} */,
  {32'h4552a8e4, 32'h457ff964} /* (10, 3, 1) {real, imag} */,
  {32'h45b7e3a4, 32'h00000000} /* (10, 3, 0) {real, imag} */,
  {32'h455171fe, 32'hc5814cc4} /* (10, 2, 31) {real, imag} */,
  {32'h438c4717, 32'h44995146} /* (10, 2, 30) {real, imag} */,
  {32'hc2f60ed9, 32'h408cffd0} /* (10, 2, 29) {real, imag} */,
  {32'hc3273098, 32'h43b4af38} /* (10, 2, 28) {real, imag} */,
  {32'hc31053bc, 32'hc3088da5} /* (10, 2, 27) {real, imag} */,
  {32'hc2760a03, 32'h42b50860} /* (10, 2, 26) {real, imag} */,
  {32'h41ea5f7d, 32'h40de5ba8} /* (10, 2, 25) {real, imag} */,
  {32'h42543e7b, 32'h42ac5d5a} /* (10, 2, 24) {real, imag} */,
  {32'hc2b038e8, 32'hc214c231} /* (10, 2, 23) {real, imag} */,
  {32'h42f871fb, 32'hc212a883} /* (10, 2, 22) {real, imag} */,
  {32'hc18813b4, 32'h41c7d628} /* (10, 2, 21) {real, imag} */,
  {32'h418a20c8, 32'h418db71f} /* (10, 2, 20) {real, imag} */,
  {32'h4170fd0f, 32'h424489ec} /* (10, 2, 19) {real, imag} */,
  {32'h417d2be8, 32'hc1a3b33e} /* (10, 2, 18) {real, imag} */,
  {32'h4251fff7, 32'hc1e48b18} /* (10, 2, 17) {real, imag} */,
  {32'hc2c8eb42, 32'h00000000} /* (10, 2, 16) {real, imag} */,
  {32'h4251fff7, 32'h41e48b18} /* (10, 2, 15) {real, imag} */,
  {32'h417d2be8, 32'h41a3b33e} /* (10, 2, 14) {real, imag} */,
  {32'h4170fd0f, 32'hc24489ec} /* (10, 2, 13) {real, imag} */,
  {32'h418a20c8, 32'hc18db71f} /* (10, 2, 12) {real, imag} */,
  {32'hc18813b4, 32'hc1c7d628} /* (10, 2, 11) {real, imag} */,
  {32'h42f871fb, 32'h4212a883} /* (10, 2, 10) {real, imag} */,
  {32'hc2b038e8, 32'h4214c231} /* (10, 2, 9) {real, imag} */,
  {32'h42543e7b, 32'hc2ac5d5a} /* (10, 2, 8) {real, imag} */,
  {32'h41ea5f7d, 32'hc0de5ba8} /* (10, 2, 7) {real, imag} */,
  {32'hc2760a03, 32'hc2b50860} /* (10, 2, 6) {real, imag} */,
  {32'hc31053bc, 32'h43088da5} /* (10, 2, 5) {real, imag} */,
  {32'hc3273098, 32'hc3b4af38} /* (10, 2, 4) {real, imag} */,
  {32'hc2f60ed9, 32'hc08cffd0} /* (10, 2, 3) {real, imag} */,
  {32'h438c4717, 32'hc4995146} /* (10, 2, 2) {real, imag} */,
  {32'h455171fe, 32'h45814cc4} /* (10, 2, 1) {real, imag} */,
  {32'h45b1a273, 32'h00000000} /* (10, 2, 0) {real, imag} */,
  {32'h455cce8c, 32'hc5700414} /* (10, 1, 31) {real, imag} */,
  {32'h4258e1b0, 32'h44840658} /* (10, 1, 30) {real, imag} */,
  {32'hc364d818, 32'hc315a417} /* (10, 1, 29) {real, imag} */,
  {32'hc2a1dc1b, 32'h43bd4f8c} /* (10, 1, 28) {real, imag} */,
  {32'hc3452764, 32'hc27d14a6} /* (10, 1, 27) {real, imag} */,
  {32'hc2957245, 32'h42661a22} /* (10, 1, 26) {real, imag} */,
  {32'h4200e6a7, 32'h411f12f8} /* (10, 1, 25) {real, imag} */,
  {32'h42896a7f, 32'h418d7caa} /* (10, 1, 24) {real, imag} */,
  {32'h4194fc92, 32'h42403ac6} /* (10, 1, 23) {real, imag} */,
  {32'hc296106b, 32'hc0fe4d47} /* (10, 1, 22) {real, imag} */,
  {32'h4243964d, 32'hc1ad895a} /* (10, 1, 21) {real, imag} */,
  {32'h40f33b10, 32'h424cf6f5} /* (10, 1, 20) {real, imag} */,
  {32'hc2801d03, 32'hc2378c60} /* (10, 1, 19) {real, imag} */,
  {32'h416f8404, 32'h4120e584} /* (10, 1, 18) {real, imag} */,
  {32'hc214a176, 32'h41b40798} /* (10, 1, 17) {real, imag} */,
  {32'hc0cd6ab7, 32'h00000000} /* (10, 1, 16) {real, imag} */,
  {32'hc214a176, 32'hc1b40798} /* (10, 1, 15) {real, imag} */,
  {32'h416f8404, 32'hc120e584} /* (10, 1, 14) {real, imag} */,
  {32'hc2801d03, 32'h42378c60} /* (10, 1, 13) {real, imag} */,
  {32'h40f33b10, 32'hc24cf6f5} /* (10, 1, 12) {real, imag} */,
  {32'h4243964d, 32'h41ad895a} /* (10, 1, 11) {real, imag} */,
  {32'hc296106b, 32'h40fe4d47} /* (10, 1, 10) {real, imag} */,
  {32'h4194fc92, 32'hc2403ac6} /* (10, 1, 9) {real, imag} */,
  {32'h42896a7f, 32'hc18d7caa} /* (10, 1, 8) {real, imag} */,
  {32'h4200e6a7, 32'hc11f12f8} /* (10, 1, 7) {real, imag} */,
  {32'hc2957245, 32'hc2661a22} /* (10, 1, 6) {real, imag} */,
  {32'hc3452764, 32'h427d14a6} /* (10, 1, 5) {real, imag} */,
  {32'hc2a1dc1b, 32'hc3bd4f8c} /* (10, 1, 4) {real, imag} */,
  {32'hc364d818, 32'h4315a417} /* (10, 1, 3) {real, imag} */,
  {32'h4258e1b0, 32'hc4840658} /* (10, 1, 2) {real, imag} */,
  {32'h455cce8c, 32'h45700414} /* (10, 1, 1) {real, imag} */,
  {32'h45b13a39, 32'h00000000} /* (10, 1, 0) {real, imag} */,
  {32'h456692e7, 32'hc5409ce6} /* (10, 0, 31) {real, imag} */,
  {32'hc36298f4, 32'h443ae223} /* (10, 0, 30) {real, imag} */,
  {32'hc325de0a, 32'hc24480a1} /* (10, 0, 29) {real, imag} */,
  {32'hc25855e4, 32'h43764c32} /* (10, 0, 28) {real, imag} */,
  {32'hc342ec62, 32'hc1aa8060} /* (10, 0, 27) {real, imag} */,
  {32'h3e855a00, 32'h414067d0} /* (10, 0, 26) {real, imag} */,
  {32'h4262f2d6, 32'hc15cc855} /* (10, 0, 25) {real, imag} */,
  {32'h408fe5a0, 32'hc1b21fcc} /* (10, 0, 24) {real, imag} */,
  {32'h41873a0a, 32'hbfcb3510} /* (10, 0, 23) {real, imag} */,
  {32'hc284730e, 32'hc139438a} /* (10, 0, 22) {real, imag} */,
  {32'h41ccd6f4, 32'h422358e5} /* (10, 0, 21) {real, imag} */,
  {32'hc10c10e8, 32'hc198a098} /* (10, 0, 20) {real, imag} */,
  {32'h423cc8c2, 32'hc10df9ed} /* (10, 0, 19) {real, imag} */,
  {32'hc0ef85b0, 32'h41d3c590} /* (10, 0, 18) {real, imag} */,
  {32'hc219ab63, 32'h3f560c00} /* (10, 0, 17) {real, imag} */,
  {32'h4162e64c, 32'h00000000} /* (10, 0, 16) {real, imag} */,
  {32'hc219ab63, 32'hbf560c00} /* (10, 0, 15) {real, imag} */,
  {32'hc0ef85b0, 32'hc1d3c590} /* (10, 0, 14) {real, imag} */,
  {32'h423cc8c2, 32'h410df9ed} /* (10, 0, 13) {real, imag} */,
  {32'hc10c10e8, 32'h4198a098} /* (10, 0, 12) {real, imag} */,
  {32'h41ccd6f4, 32'hc22358e5} /* (10, 0, 11) {real, imag} */,
  {32'hc284730e, 32'h4139438a} /* (10, 0, 10) {real, imag} */,
  {32'h41873a0a, 32'h3fcb3510} /* (10, 0, 9) {real, imag} */,
  {32'h408fe5a0, 32'h41b21fcc} /* (10, 0, 8) {real, imag} */,
  {32'h4262f2d6, 32'h415cc855} /* (10, 0, 7) {real, imag} */,
  {32'h3e855a00, 32'hc14067d0} /* (10, 0, 6) {real, imag} */,
  {32'hc342ec62, 32'h41aa8060} /* (10, 0, 5) {real, imag} */,
  {32'hc25855e4, 32'hc3764c32} /* (10, 0, 4) {real, imag} */,
  {32'hc325de0a, 32'h424480a1} /* (10, 0, 3) {real, imag} */,
  {32'hc36298f4, 32'hc43ae223} /* (10, 0, 2) {real, imag} */,
  {32'h456692e7, 32'h45409ce6} /* (10, 0, 1) {real, imag} */,
  {32'h45b1008c, 32'h00000000} /* (10, 0, 0) {real, imag} */,
  {32'h457763e7, 32'hc5116a1f} /* (9, 31, 31) {real, imag} */,
  {32'hc455096a, 32'h4436d006} /* (9, 31, 30) {real, imag} */,
  {32'hc2366328, 32'hc2c3517e} /* (9, 31, 29) {real, imag} */,
  {32'h42ff1a90, 32'h42cc7c04} /* (9, 31, 28) {real, imag} */,
  {32'hc32f353b, 32'hc102c3c8} /* (9, 31, 27) {real, imag} */,
  {32'h420c2070, 32'h42077a6c} /* (9, 31, 26) {real, imag} */,
  {32'hc2086744, 32'h4178b916} /* (9, 31, 25) {real, imag} */,
  {32'hc225c60c, 32'hbfd358c0} /* (9, 31, 24) {real, imag} */,
  {32'h428b0064, 32'h41ae2c48} /* (9, 31, 23) {real, imag} */,
  {32'hc16e2b1c, 32'h408e2ab6} /* (9, 31, 22) {real, imag} */,
  {32'h41e1e30a, 32'hc19bc81e} /* (9, 31, 21) {real, imag} */,
  {32'h4274afa6, 32'hc234cbe5} /* (9, 31, 20) {real, imag} */,
  {32'h413faac0, 32'hc1b9bc2e} /* (9, 31, 19) {real, imag} */,
  {32'hc24dac79, 32'hc14e3608} /* (9, 31, 18) {real, imag} */,
  {32'h3fbb02d4, 32'h40bd23f0} /* (9, 31, 17) {real, imag} */,
  {32'hc0c1b1bc, 32'h00000000} /* (9, 31, 16) {real, imag} */,
  {32'h3fbb02d4, 32'hc0bd23f0} /* (9, 31, 15) {real, imag} */,
  {32'hc24dac79, 32'h414e3608} /* (9, 31, 14) {real, imag} */,
  {32'h413faac0, 32'h41b9bc2e} /* (9, 31, 13) {real, imag} */,
  {32'h4274afa6, 32'h4234cbe5} /* (9, 31, 12) {real, imag} */,
  {32'h41e1e30a, 32'h419bc81e} /* (9, 31, 11) {real, imag} */,
  {32'hc16e2b1c, 32'hc08e2ab6} /* (9, 31, 10) {real, imag} */,
  {32'h428b0064, 32'hc1ae2c48} /* (9, 31, 9) {real, imag} */,
  {32'hc225c60c, 32'h3fd358c0} /* (9, 31, 8) {real, imag} */,
  {32'hc2086744, 32'hc178b916} /* (9, 31, 7) {real, imag} */,
  {32'h420c2070, 32'hc2077a6c} /* (9, 31, 6) {real, imag} */,
  {32'hc32f353b, 32'h4102c3c8} /* (9, 31, 5) {real, imag} */,
  {32'h42ff1a90, 32'hc2cc7c04} /* (9, 31, 4) {real, imag} */,
  {32'hc2366328, 32'h42c3517e} /* (9, 31, 3) {real, imag} */,
  {32'hc455096a, 32'hc436d006} /* (9, 31, 2) {real, imag} */,
  {32'h457763e7, 32'h45116a1f} /* (9, 31, 1) {real, imag} */,
  {32'h45af322b, 32'h00000000} /* (9, 31, 0) {real, imag} */,
  {32'h458ee383, 32'hc4e757d4} /* (9, 30, 31) {real, imag} */,
  {32'hc495d64e, 32'h441d7709} /* (9, 30, 30) {real, imag} */,
  {32'hc205e090, 32'hc2b42c85} /* (9, 30, 29) {real, imag} */,
  {32'h4319839a, 32'h421a30d0} /* (9, 30, 28) {real, imag} */,
  {32'hc3697fbd, 32'h416e3358} /* (9, 30, 27) {real, imag} */,
  {32'h4219a3cd, 32'hc1cc8213} /* (9, 30, 26) {real, imag} */,
  {32'h424a027e, 32'h427d5495} /* (9, 30, 25) {real, imag} */,
  {32'hc22b06f6, 32'hc0a3e1a0} /* (9, 30, 24) {real, imag} */,
  {32'h42e9e25b, 32'h4111f938} /* (9, 30, 23) {real, imag} */,
  {32'h41d2cf8c, 32'h43018678} /* (9, 30, 22) {real, imag} */,
  {32'hc085d998, 32'h42c1d71a} /* (9, 30, 21) {real, imag} */,
  {32'h430017da, 32'hc210619a} /* (9, 30, 20) {real, imag} */,
  {32'h42bdac41, 32'hc2f833d2} /* (9, 30, 19) {real, imag} */,
  {32'h412e4dec, 32'h41fd1200} /* (9, 30, 18) {real, imag} */,
  {32'hc1a47567, 32'hc086d428} /* (9, 30, 17) {real, imag} */,
  {32'hc19eca90, 32'h00000000} /* (9, 30, 16) {real, imag} */,
  {32'hc1a47567, 32'h4086d428} /* (9, 30, 15) {real, imag} */,
  {32'h412e4dec, 32'hc1fd1200} /* (9, 30, 14) {real, imag} */,
  {32'h42bdac41, 32'h42f833d2} /* (9, 30, 13) {real, imag} */,
  {32'h430017da, 32'h4210619a} /* (9, 30, 12) {real, imag} */,
  {32'hc085d998, 32'hc2c1d71a} /* (9, 30, 11) {real, imag} */,
  {32'h41d2cf8c, 32'hc3018678} /* (9, 30, 10) {real, imag} */,
  {32'h42e9e25b, 32'hc111f938} /* (9, 30, 9) {real, imag} */,
  {32'hc22b06f6, 32'h40a3e1a0} /* (9, 30, 8) {real, imag} */,
  {32'h424a027e, 32'hc27d5495} /* (9, 30, 7) {real, imag} */,
  {32'h4219a3cd, 32'h41cc8213} /* (9, 30, 6) {real, imag} */,
  {32'hc3697fbd, 32'hc16e3358} /* (9, 30, 5) {real, imag} */,
  {32'h4319839a, 32'hc21a30d0} /* (9, 30, 4) {real, imag} */,
  {32'hc205e090, 32'h42b42c85} /* (9, 30, 3) {real, imag} */,
  {32'hc495d64e, 32'hc41d7709} /* (9, 30, 2) {real, imag} */,
  {32'h458ee383, 32'h44e757d4} /* (9, 30, 1) {real, imag} */,
  {32'h45b45a47, 32'h00000000} /* (9, 30, 0) {real, imag} */,
  {32'h459968cd, 32'hc4c09a44} /* (9, 29, 31) {real, imag} */,
  {32'hc4adfaf9, 32'h441d52bc} /* (9, 29, 30) {real, imag} */,
  {32'h4218c36a, 32'hc288ac1f} /* (9, 29, 29) {real, imag} */,
  {32'h425933d7, 32'h410119d0} /* (9, 29, 28) {real, imag} */,
  {32'hc34012a4, 32'hc28ee97f} /* (9, 29, 27) {real, imag} */,
  {32'hc2a88e80, 32'hc00ac0f0} /* (9, 29, 26) {real, imag} */,
  {32'hc27975ee, 32'hc312c82e} /* (9, 29, 25) {real, imag} */,
  {32'hc1f2e1ea, 32'h42102df0} /* (9, 29, 24) {real, imag} */,
  {32'h42314df1, 32'hc28972ca} /* (9, 29, 23) {real, imag} */,
  {32'hc208806a, 32'h427c3bfc} /* (9, 29, 22) {real, imag} */,
  {32'hc2932c0e, 32'h3f861d10} /* (9, 29, 21) {real, imag} */,
  {32'hc0af3f74, 32'h42d91383} /* (9, 29, 20) {real, imag} */,
  {32'hc2af8d86, 32'h411bedd8} /* (9, 29, 19) {real, imag} */,
  {32'hc1c43059, 32'h41ebe415} /* (9, 29, 18) {real, imag} */,
  {32'hc0c663a0, 32'hc1556086} /* (9, 29, 17) {real, imag} */,
  {32'hc1839f50, 32'h00000000} /* (9, 29, 16) {real, imag} */,
  {32'hc0c663a0, 32'h41556086} /* (9, 29, 15) {real, imag} */,
  {32'hc1c43059, 32'hc1ebe415} /* (9, 29, 14) {real, imag} */,
  {32'hc2af8d86, 32'hc11bedd8} /* (9, 29, 13) {real, imag} */,
  {32'hc0af3f74, 32'hc2d91383} /* (9, 29, 12) {real, imag} */,
  {32'hc2932c0e, 32'hbf861d10} /* (9, 29, 11) {real, imag} */,
  {32'hc208806a, 32'hc27c3bfc} /* (9, 29, 10) {real, imag} */,
  {32'h42314df1, 32'h428972ca} /* (9, 29, 9) {real, imag} */,
  {32'hc1f2e1ea, 32'hc2102df0} /* (9, 29, 8) {real, imag} */,
  {32'hc27975ee, 32'h4312c82e} /* (9, 29, 7) {real, imag} */,
  {32'hc2a88e80, 32'h400ac0f0} /* (9, 29, 6) {real, imag} */,
  {32'hc34012a4, 32'h428ee97f} /* (9, 29, 5) {real, imag} */,
  {32'h425933d7, 32'hc10119d0} /* (9, 29, 4) {real, imag} */,
  {32'h4218c36a, 32'h4288ac1f} /* (9, 29, 3) {real, imag} */,
  {32'hc4adfaf9, 32'hc41d52bc} /* (9, 29, 2) {real, imag} */,
  {32'h459968cd, 32'h44c09a44} /* (9, 29, 1) {real, imag} */,
  {32'h45b1f1cf, 32'h00000000} /* (9, 29, 0) {real, imag} */,
  {32'h45a1369f, 32'hc48fbcb2} /* (9, 28, 31) {real, imag} */,
  {32'hc4cd74c0, 32'h4410dcb1} /* (9, 28, 30) {real, imag} */,
  {32'h431f7faa, 32'h4153508c} /* (9, 28, 29) {real, imag} */,
  {32'h434366e6, 32'hc2a5470c} /* (9, 28, 28) {real, imag} */,
  {32'hc381f52b, 32'hc293200f} /* (9, 28, 27) {real, imag} */,
  {32'hc2d6e7a6, 32'hc2334e60} /* (9, 28, 26) {real, imag} */,
  {32'h42dbbdf6, 32'hc31c555c} /* (9, 28, 25) {real, imag} */,
  {32'hc1aee018, 32'h41b42caa} /* (9, 28, 24) {real, imag} */,
  {32'hc2acad8a, 32'hc2d76151} /* (9, 28, 23) {real, imag} */,
  {32'h3f4d73f0, 32'h4192bc0e} /* (9, 28, 22) {real, imag} */,
  {32'hc2acda0e, 32'h4287ddc2} /* (9, 28, 21) {real, imag} */,
  {32'h41b4b1d4, 32'h4222e449} /* (9, 28, 20) {real, imag} */,
  {32'h4292801a, 32'h41fafbb8} /* (9, 28, 19) {real, imag} */,
  {32'hc285bc66, 32'h424739f4} /* (9, 28, 18) {real, imag} */,
  {32'hc307991f, 32'h42444e21} /* (9, 28, 17) {real, imag} */,
  {32'h42abfa5d, 32'h00000000} /* (9, 28, 16) {real, imag} */,
  {32'hc307991f, 32'hc2444e21} /* (9, 28, 15) {real, imag} */,
  {32'hc285bc66, 32'hc24739f4} /* (9, 28, 14) {real, imag} */,
  {32'h4292801a, 32'hc1fafbb8} /* (9, 28, 13) {real, imag} */,
  {32'h41b4b1d4, 32'hc222e449} /* (9, 28, 12) {real, imag} */,
  {32'hc2acda0e, 32'hc287ddc2} /* (9, 28, 11) {real, imag} */,
  {32'h3f4d73f0, 32'hc192bc0e} /* (9, 28, 10) {real, imag} */,
  {32'hc2acad8a, 32'h42d76151} /* (9, 28, 9) {real, imag} */,
  {32'hc1aee018, 32'hc1b42caa} /* (9, 28, 8) {real, imag} */,
  {32'h42dbbdf6, 32'h431c555c} /* (9, 28, 7) {real, imag} */,
  {32'hc2d6e7a6, 32'h42334e60} /* (9, 28, 6) {real, imag} */,
  {32'hc381f52b, 32'h4293200f} /* (9, 28, 5) {real, imag} */,
  {32'h434366e6, 32'h42a5470c} /* (9, 28, 4) {real, imag} */,
  {32'h431f7faa, 32'hc153508c} /* (9, 28, 3) {real, imag} */,
  {32'hc4cd74c0, 32'hc410dcb1} /* (9, 28, 2) {real, imag} */,
  {32'h45a1369f, 32'h448fbcb2} /* (9, 28, 1) {real, imag} */,
  {32'h45b10cf8, 32'h00000000} /* (9, 28, 0) {real, imag} */,
  {32'h45a41d81, 32'hc457b88e} /* (9, 27, 31) {real, imag} */,
  {32'hc4e03bd8, 32'h43e6f0a2} /* (9, 27, 30) {real, imag} */,
  {32'hc3025fbf, 32'h42c37b06} /* (9, 27, 29) {real, imag} */,
  {32'h439b2bf3, 32'hc25268b0} /* (9, 27, 28) {real, imag} */,
  {32'hc2829226, 32'hc2309c5c} /* (9, 27, 27) {real, imag} */,
  {32'hc2f755c0, 32'hc0b0d660} /* (9, 27, 26) {real, imag} */,
  {32'h4271d62b, 32'hc1b1ee84} /* (9, 27, 25) {real, imag} */,
  {32'hc2ab39ea, 32'h42bb994a} /* (9, 27, 24) {real, imag} */,
  {32'h429d6f93, 32'h422113e3} /* (9, 27, 23) {real, imag} */,
  {32'h41be71c6, 32'hbf296020} /* (9, 27, 22) {real, imag} */,
  {32'hc29a33bd, 32'h415a8c14} /* (9, 27, 21) {real, imag} */,
  {32'hc2169538, 32'h42452436} /* (9, 27, 20) {real, imag} */,
  {32'h42d27e9e, 32'hc1e594a0} /* (9, 27, 19) {real, imag} */,
  {32'h427145f8, 32'h427d0457} /* (9, 27, 18) {real, imag} */,
  {32'hc265baa3, 32'hc2952f57} /* (9, 27, 17) {real, imag} */,
  {32'hc2cbec3a, 32'h00000000} /* (9, 27, 16) {real, imag} */,
  {32'hc265baa3, 32'h42952f57} /* (9, 27, 15) {real, imag} */,
  {32'h427145f8, 32'hc27d0457} /* (9, 27, 14) {real, imag} */,
  {32'h42d27e9e, 32'h41e594a0} /* (9, 27, 13) {real, imag} */,
  {32'hc2169538, 32'hc2452436} /* (9, 27, 12) {real, imag} */,
  {32'hc29a33bd, 32'hc15a8c14} /* (9, 27, 11) {real, imag} */,
  {32'h41be71c6, 32'h3f296020} /* (9, 27, 10) {real, imag} */,
  {32'h429d6f93, 32'hc22113e3} /* (9, 27, 9) {real, imag} */,
  {32'hc2ab39ea, 32'hc2bb994a} /* (9, 27, 8) {real, imag} */,
  {32'h4271d62b, 32'h41b1ee84} /* (9, 27, 7) {real, imag} */,
  {32'hc2f755c0, 32'h40b0d660} /* (9, 27, 6) {real, imag} */,
  {32'hc2829226, 32'h42309c5c} /* (9, 27, 5) {real, imag} */,
  {32'h439b2bf3, 32'h425268b0} /* (9, 27, 4) {real, imag} */,
  {32'hc3025fbf, 32'hc2c37b06} /* (9, 27, 3) {real, imag} */,
  {32'hc4e03bd8, 32'hc3e6f0a2} /* (9, 27, 2) {real, imag} */,
  {32'h45a41d81, 32'h4457b88e} /* (9, 27, 1) {real, imag} */,
  {32'h45adc4a0, 32'h00000000} /* (9, 27, 0) {real, imag} */,
  {32'h459f97e5, 32'hc4241b26} /* (9, 26, 31) {real, imag} */,
  {32'hc4dde798, 32'h4384580c} /* (9, 26, 30) {real, imag} */,
  {32'hc213bf30, 32'h42950740} /* (9, 26, 29) {real, imag} */,
  {32'h434a411a, 32'hc293511e} /* (9, 26, 28) {real, imag} */,
  {32'hc32882d4, 32'h41e880cf} /* (9, 26, 27) {real, imag} */,
  {32'hc280cde0, 32'h41533bf8} /* (9, 26, 26) {real, imag} */,
  {32'hc22672aa, 32'h40cbcde0} /* (9, 26, 25) {real, imag} */,
  {32'hc188d24c, 32'h43482412} /* (9, 26, 24) {real, imag} */,
  {32'h42f35db3, 32'h4012eb84} /* (9, 26, 23) {real, imag} */,
  {32'hc26689ba, 32'hc23bc230} /* (9, 26, 22) {real, imag} */,
  {32'h42826c1d, 32'h41f7fcca} /* (9, 26, 21) {real, imag} */,
  {32'h4118b95f, 32'hc04f6988} /* (9, 26, 20) {real, imag} */,
  {32'hc2b3296c, 32'hc2022b14} /* (9, 26, 19) {real, imag} */,
  {32'hc22481e2, 32'hc0a5c2b0} /* (9, 26, 18) {real, imag} */,
  {32'h41c5f9ba, 32'h41d0e777} /* (9, 26, 17) {real, imag} */,
  {32'h41c97b48, 32'h00000000} /* (9, 26, 16) {real, imag} */,
  {32'h41c5f9ba, 32'hc1d0e777} /* (9, 26, 15) {real, imag} */,
  {32'hc22481e2, 32'h40a5c2b0} /* (9, 26, 14) {real, imag} */,
  {32'hc2b3296c, 32'h42022b14} /* (9, 26, 13) {real, imag} */,
  {32'h4118b95f, 32'h404f6988} /* (9, 26, 12) {real, imag} */,
  {32'h42826c1d, 32'hc1f7fcca} /* (9, 26, 11) {real, imag} */,
  {32'hc26689ba, 32'h423bc230} /* (9, 26, 10) {real, imag} */,
  {32'h42f35db3, 32'hc012eb84} /* (9, 26, 9) {real, imag} */,
  {32'hc188d24c, 32'hc3482412} /* (9, 26, 8) {real, imag} */,
  {32'hc22672aa, 32'hc0cbcde0} /* (9, 26, 7) {real, imag} */,
  {32'hc280cde0, 32'hc1533bf8} /* (9, 26, 6) {real, imag} */,
  {32'hc32882d4, 32'hc1e880cf} /* (9, 26, 5) {real, imag} */,
  {32'h434a411a, 32'h4293511e} /* (9, 26, 4) {real, imag} */,
  {32'hc213bf30, 32'hc2950740} /* (9, 26, 3) {real, imag} */,
  {32'hc4dde798, 32'hc384580c} /* (9, 26, 2) {real, imag} */,
  {32'h459f97e5, 32'h44241b26} /* (9, 26, 1) {real, imag} */,
  {32'h45a84759, 32'h00000000} /* (9, 26, 0) {real, imag} */,
  {32'h45972706, 32'hc3baa238} /* (9, 25, 31) {real, imag} */,
  {32'hc4cd72f3, 32'h43873dee} /* (9, 25, 30) {real, imag} */,
  {32'hc2ab52b6, 32'h408612f0} /* (9, 25, 29) {real, imag} */,
  {32'h42b33a65, 32'hc2d9be1e} /* (9, 25, 28) {real, imag} */,
  {32'hc3505bf4, 32'h4283abfd} /* (9, 25, 27) {real, imag} */,
  {32'hc2208c60, 32'hc2278e86} /* (9, 25, 26) {real, imag} */,
  {32'h4282e64c, 32'h42d8c89c} /* (9, 25, 25) {real, imag} */,
  {32'h42711a3e, 32'h430ad227} /* (9, 25, 24) {real, imag} */,
  {32'h3f449660, 32'hc16fb2ee} /* (9, 25, 23) {real, imag} */,
  {32'h4263798f, 32'hc3252f08} /* (9, 25, 22) {real, imag} */,
  {32'h41ff5294, 32'h42750308} /* (9, 25, 21) {real, imag} */,
  {32'hc2933757, 32'h41c8e554} /* (9, 25, 20) {real, imag} */,
  {32'hc2a3e279, 32'hc12626ad} /* (9, 25, 19) {real, imag} */,
  {32'h41c00fe2, 32'h430214ae} /* (9, 25, 18) {real, imag} */,
  {32'h408f286a, 32'h4157f966} /* (9, 25, 17) {real, imag} */,
  {32'h41a56edd, 32'h00000000} /* (9, 25, 16) {real, imag} */,
  {32'h408f286a, 32'hc157f966} /* (9, 25, 15) {real, imag} */,
  {32'h41c00fe2, 32'hc30214ae} /* (9, 25, 14) {real, imag} */,
  {32'hc2a3e279, 32'h412626ad} /* (9, 25, 13) {real, imag} */,
  {32'hc2933757, 32'hc1c8e554} /* (9, 25, 12) {real, imag} */,
  {32'h41ff5294, 32'hc2750308} /* (9, 25, 11) {real, imag} */,
  {32'h4263798f, 32'h43252f08} /* (9, 25, 10) {real, imag} */,
  {32'h3f449660, 32'h416fb2ee} /* (9, 25, 9) {real, imag} */,
  {32'h42711a3e, 32'hc30ad227} /* (9, 25, 8) {real, imag} */,
  {32'h4282e64c, 32'hc2d8c89c} /* (9, 25, 7) {real, imag} */,
  {32'hc2208c60, 32'h42278e86} /* (9, 25, 6) {real, imag} */,
  {32'hc3505bf4, 32'hc283abfd} /* (9, 25, 5) {real, imag} */,
  {32'h42b33a65, 32'h42d9be1e} /* (9, 25, 4) {real, imag} */,
  {32'hc2ab52b6, 32'hc08612f0} /* (9, 25, 3) {real, imag} */,
  {32'hc4cd72f3, 32'hc3873dee} /* (9, 25, 2) {real, imag} */,
  {32'h45972706, 32'h43baa238} /* (9, 25, 1) {real, imag} */,
  {32'h459c3cd4, 32'h00000000} /* (9, 25, 0) {real, imag} */,
  {32'h45818981, 32'hc31f48e8} /* (9, 24, 31) {real, imag} */,
  {32'hc4b22063, 32'h439adee7} /* (9, 24, 30) {real, imag} */,
  {32'hc343110e, 32'hc306fed8} /* (9, 24, 29) {real, imag} */,
  {32'h43967d17, 32'h412806e0} /* (9, 24, 28) {real, imag} */,
  {32'hc3637fe7, 32'hc1b27bfd} /* (9, 24, 27) {real, imag} */,
  {32'hc2a72041, 32'hc2b0c35b} /* (9, 24, 26) {real, imag} */,
  {32'h425f916a, 32'hc2b0f486} /* (9, 24, 25) {real, imag} */,
  {32'hc34d5843, 32'h4326df2b} /* (9, 24, 24) {real, imag} */,
  {32'hc209d3fe, 32'hc3096206} /* (9, 24, 23) {real, imag} */,
  {32'h3f493da0, 32'h42e47727} /* (9, 24, 22) {real, imag} */,
  {32'hc2ae5ce6, 32'h42426866} /* (9, 24, 21) {real, imag} */,
  {32'h415f1028, 32'hc1a9b786} /* (9, 24, 20) {real, imag} */,
  {32'h4248fb5a, 32'h41b60c2d} /* (9, 24, 19) {real, imag} */,
  {32'h42174c28, 32'h42d7949b} /* (9, 24, 18) {real, imag} */,
  {32'h41eff92e, 32'hc1d1c60c} /* (9, 24, 17) {real, imag} */,
  {32'h420a79ac, 32'h00000000} /* (9, 24, 16) {real, imag} */,
  {32'h41eff92e, 32'h41d1c60c} /* (9, 24, 15) {real, imag} */,
  {32'h42174c28, 32'hc2d7949b} /* (9, 24, 14) {real, imag} */,
  {32'h4248fb5a, 32'hc1b60c2d} /* (9, 24, 13) {real, imag} */,
  {32'h415f1028, 32'h41a9b786} /* (9, 24, 12) {real, imag} */,
  {32'hc2ae5ce6, 32'hc2426866} /* (9, 24, 11) {real, imag} */,
  {32'h3f493da0, 32'hc2e47727} /* (9, 24, 10) {real, imag} */,
  {32'hc209d3fe, 32'h43096206} /* (9, 24, 9) {real, imag} */,
  {32'hc34d5843, 32'hc326df2b} /* (9, 24, 8) {real, imag} */,
  {32'h425f916a, 32'h42b0f486} /* (9, 24, 7) {real, imag} */,
  {32'hc2a72041, 32'h42b0c35b} /* (9, 24, 6) {real, imag} */,
  {32'hc3637fe7, 32'h41b27bfd} /* (9, 24, 5) {real, imag} */,
  {32'h43967d17, 32'hc12806e0} /* (9, 24, 4) {real, imag} */,
  {32'hc343110e, 32'h4306fed8} /* (9, 24, 3) {real, imag} */,
  {32'hc4b22063, 32'hc39adee7} /* (9, 24, 2) {real, imag} */,
  {32'h45818981, 32'h431f48e8} /* (9, 24, 1) {real, imag} */,
  {32'h4584cf5a, 32'h00000000} /* (9, 24, 0) {real, imag} */,
  {32'h454e33da, 32'hc333120c} /* (9, 23, 31) {real, imag} */,
  {32'hc49b486b, 32'h4372c863} /* (9, 23, 30) {real, imag} */,
  {32'hc2f17542, 32'hc1c5f0eb} /* (9, 23, 29) {real, imag} */,
  {32'h43804937, 32'hc2d63244} /* (9, 23, 28) {real, imag} */,
  {32'hc3750eaa, 32'h42ffd0be} /* (9, 23, 27) {real, imag} */,
  {32'hc22606a8, 32'h42648624} /* (9, 23, 26) {real, imag} */,
  {32'h42a153b9, 32'hc2420dd8} /* (9, 23, 25) {real, imag} */,
  {32'h3ed11bc0, 32'h40b342a8} /* (9, 23, 24) {real, imag} */,
  {32'hc267e4d5, 32'hc2077cf7} /* (9, 23, 23) {real, imag} */,
  {32'h4139f7db, 32'h429d0b4d} /* (9, 23, 22) {real, imag} */,
  {32'h413cc99c, 32'h4287759c} /* (9, 23, 21) {real, imag} */,
  {32'hc2492794, 32'hc288176e} /* (9, 23, 20) {real, imag} */,
  {32'hc0d95d72, 32'h424de485} /* (9, 23, 19) {real, imag} */,
  {32'hc215b147, 32'h42022e40} /* (9, 23, 18) {real, imag} */,
  {32'hc223988b, 32'hc2bc1242} /* (9, 23, 17) {real, imag} */,
  {32'h426ac61e, 32'h00000000} /* (9, 23, 16) {real, imag} */,
  {32'hc223988b, 32'h42bc1242} /* (9, 23, 15) {real, imag} */,
  {32'hc215b147, 32'hc2022e40} /* (9, 23, 14) {real, imag} */,
  {32'hc0d95d72, 32'hc24de485} /* (9, 23, 13) {real, imag} */,
  {32'hc2492794, 32'h4288176e} /* (9, 23, 12) {real, imag} */,
  {32'h413cc99c, 32'hc287759c} /* (9, 23, 11) {real, imag} */,
  {32'h4139f7db, 32'hc29d0b4d} /* (9, 23, 10) {real, imag} */,
  {32'hc267e4d5, 32'h42077cf7} /* (9, 23, 9) {real, imag} */,
  {32'h3ed11bc0, 32'hc0b342a8} /* (9, 23, 8) {real, imag} */,
  {32'h42a153b9, 32'h42420dd8} /* (9, 23, 7) {real, imag} */,
  {32'hc22606a8, 32'hc2648624} /* (9, 23, 6) {real, imag} */,
  {32'hc3750eaa, 32'hc2ffd0be} /* (9, 23, 5) {real, imag} */,
  {32'h43804937, 32'h42d63244} /* (9, 23, 4) {real, imag} */,
  {32'hc2f17542, 32'h41c5f0eb} /* (9, 23, 3) {real, imag} */,
  {32'hc49b486b, 32'hc372c863} /* (9, 23, 2) {real, imag} */,
  {32'h454e33da, 32'h4333120c} /* (9, 23, 1) {real, imag} */,
  {32'h455373fe, 32'h00000000} /* (9, 23, 0) {real, imag} */,
  {32'h450f0cd4, 32'hc346abc6} /* (9, 22, 31) {real, imag} */,
  {32'hc455ae5c, 32'h42996730} /* (9, 22, 30) {real, imag} */,
  {32'hc272bedc, 32'h430928ae} /* (9, 22, 29) {real, imag} */,
  {32'h42775afe, 32'hc2c0e412} /* (9, 22, 28) {real, imag} */,
  {32'hc3a2912c, 32'h4266bce4} /* (9, 22, 27) {real, imag} */,
  {32'hc21e9fd0, 32'h41932362} /* (9, 22, 26) {real, imag} */,
  {32'hc2afa2fb, 32'h42aaacea} /* (9, 22, 25) {real, imag} */,
  {32'hc1b306dc, 32'h41eff042} /* (9, 22, 24) {real, imag} */,
  {32'hc26a7d4a, 32'h422e5e20} /* (9, 22, 23) {real, imag} */,
  {32'h428df493, 32'hc1f3be1d} /* (9, 22, 22) {real, imag} */,
  {32'h4113c540, 32'hc281c8ce} /* (9, 22, 21) {real, imag} */,
  {32'h416d16c7, 32'hc1a6af21} /* (9, 22, 20) {real, imag} */,
  {32'hc20d7c51, 32'h3fab7b80} /* (9, 22, 19) {real, imag} */,
  {32'h4085e844, 32'h42795df4} /* (9, 22, 18) {real, imag} */,
  {32'h429afd2f, 32'hc2242ef2} /* (9, 22, 17) {real, imag} */,
  {32'hc2b6cb15, 32'h00000000} /* (9, 22, 16) {real, imag} */,
  {32'h429afd2f, 32'h42242ef2} /* (9, 22, 15) {real, imag} */,
  {32'h4085e844, 32'hc2795df4} /* (9, 22, 14) {real, imag} */,
  {32'hc20d7c51, 32'hbfab7b80} /* (9, 22, 13) {real, imag} */,
  {32'h416d16c7, 32'h41a6af21} /* (9, 22, 12) {real, imag} */,
  {32'h4113c540, 32'h4281c8ce} /* (9, 22, 11) {real, imag} */,
  {32'h428df493, 32'h41f3be1d} /* (9, 22, 10) {real, imag} */,
  {32'hc26a7d4a, 32'hc22e5e20} /* (9, 22, 9) {real, imag} */,
  {32'hc1b306dc, 32'hc1eff042} /* (9, 22, 8) {real, imag} */,
  {32'hc2afa2fb, 32'hc2aaacea} /* (9, 22, 7) {real, imag} */,
  {32'hc21e9fd0, 32'hc1932362} /* (9, 22, 6) {real, imag} */,
  {32'hc3a2912c, 32'hc266bce4} /* (9, 22, 5) {real, imag} */,
  {32'h42775afe, 32'h42c0e412} /* (9, 22, 4) {real, imag} */,
  {32'hc272bedc, 32'hc30928ae} /* (9, 22, 3) {real, imag} */,
  {32'hc455ae5c, 32'hc2996730} /* (9, 22, 2) {real, imag} */,
  {32'h450f0cd4, 32'h4346abc6} /* (9, 22, 1) {real, imag} */,
  {32'h451baa7e, 32'h00000000} /* (9, 22, 0) {real, imag} */,
  {32'h442276b1, 32'hc25207d8} /* (9, 21, 31) {real, imag} */,
  {32'hc36c9442, 32'hc203ed84} /* (9, 21, 30) {real, imag} */,
  {32'hc1e738eb, 32'h43443598} /* (9, 21, 29) {real, imag} */,
  {32'h42b56ee3, 32'hc184ccc4} /* (9, 21, 28) {real, imag} */,
  {32'hc314cbab, 32'h423139ed} /* (9, 21, 27) {real, imag} */,
  {32'h423ab74d, 32'hc1088f30} /* (9, 21, 26) {real, imag} */,
  {32'hc2d18561, 32'hc2ac569e} /* (9, 21, 25) {real, imag} */,
  {32'hc2bcaa7d, 32'h431cb806} /* (9, 21, 24) {real, imag} */,
  {32'hc0a7d1f0, 32'hc236f7b8} /* (9, 21, 23) {real, imag} */,
  {32'hc2328cf8, 32'hc29bc405} /* (9, 21, 22) {real, imag} */,
  {32'hc2bca0cf, 32'h422d4b51} /* (9, 21, 21) {real, imag} */,
  {32'h424849da, 32'hc310aac2} /* (9, 21, 20) {real, imag} */,
  {32'hc2830655, 32'hc2991186} /* (9, 21, 19) {real, imag} */,
  {32'h42cad2ca, 32'h42920a09} /* (9, 21, 18) {real, imag} */,
  {32'h3ffcb5f8, 32'hc2a1270e} /* (9, 21, 17) {real, imag} */,
  {32'h426c2087, 32'h00000000} /* (9, 21, 16) {real, imag} */,
  {32'h3ffcb5f8, 32'h42a1270e} /* (9, 21, 15) {real, imag} */,
  {32'h42cad2ca, 32'hc2920a09} /* (9, 21, 14) {real, imag} */,
  {32'hc2830655, 32'h42991186} /* (9, 21, 13) {real, imag} */,
  {32'h424849da, 32'h4310aac2} /* (9, 21, 12) {real, imag} */,
  {32'hc2bca0cf, 32'hc22d4b51} /* (9, 21, 11) {real, imag} */,
  {32'hc2328cf8, 32'h429bc405} /* (9, 21, 10) {real, imag} */,
  {32'hc0a7d1f0, 32'h4236f7b8} /* (9, 21, 9) {real, imag} */,
  {32'hc2bcaa7d, 32'hc31cb806} /* (9, 21, 8) {real, imag} */,
  {32'hc2d18561, 32'h42ac569e} /* (9, 21, 7) {real, imag} */,
  {32'h423ab74d, 32'h41088f30} /* (9, 21, 6) {real, imag} */,
  {32'hc314cbab, 32'hc23139ed} /* (9, 21, 5) {real, imag} */,
  {32'h42b56ee3, 32'h4184ccc4} /* (9, 21, 4) {real, imag} */,
  {32'hc1e738eb, 32'hc3443598} /* (9, 21, 3) {real, imag} */,
  {32'hc36c9442, 32'h4203ed84} /* (9, 21, 2) {real, imag} */,
  {32'h442276b1, 32'h425207d8} /* (9, 21, 1) {real, imag} */,
  {32'h448b0775, 32'h00000000} /* (9, 21, 0) {real, imag} */,
  {32'hc4a37382, 32'h42e5c240} /* (9, 20, 31) {real, imag} */,
  {32'h43fa8a88, 32'hc3772e4f} /* (9, 20, 30) {real, imag} */,
  {32'h41862aa4, 32'h4316a083} /* (9, 20, 29) {real, imag} */,
  {32'hc3316a45, 32'hc24c269c} /* (9, 20, 28) {real, imag} */,
  {32'h429fae32, 32'hc2019336} /* (9, 20, 27) {real, imag} */,
  {32'h42f8b1cc, 32'hc189f9e3} /* (9, 20, 26) {real, imag} */,
  {32'hc1a36cb9, 32'hc2185782} /* (9, 20, 25) {real, imag} */,
  {32'h4270d975, 32'hc1fe95b4} /* (9, 20, 24) {real, imag} */,
  {32'hc2b1277a, 32'hc1a1eb88} /* (9, 20, 23) {real, imag} */,
  {32'hc1bab4f0, 32'h41b4dc10} /* (9, 20, 22) {real, imag} */,
  {32'h41457a9e, 32'hc2b876e8} /* (9, 20, 21) {real, imag} */,
  {32'hc0b67292, 32'hc20135f2} /* (9, 20, 20) {real, imag} */,
  {32'h42ca447d, 32'h410c0460} /* (9, 20, 19) {real, imag} */,
  {32'h415ef817, 32'hc23ffeea} /* (9, 20, 18) {real, imag} */,
  {32'h3ea718c0, 32'h4206ff5f} /* (9, 20, 17) {real, imag} */,
  {32'h42bb0d3a, 32'h00000000} /* (9, 20, 16) {real, imag} */,
  {32'h3ea718c0, 32'hc206ff5f} /* (9, 20, 15) {real, imag} */,
  {32'h415ef817, 32'h423ffeea} /* (9, 20, 14) {real, imag} */,
  {32'h42ca447d, 32'hc10c0460} /* (9, 20, 13) {real, imag} */,
  {32'hc0b67292, 32'h420135f2} /* (9, 20, 12) {real, imag} */,
  {32'h41457a9e, 32'h42b876e8} /* (9, 20, 11) {real, imag} */,
  {32'hc1bab4f0, 32'hc1b4dc10} /* (9, 20, 10) {real, imag} */,
  {32'hc2b1277a, 32'h41a1eb88} /* (9, 20, 9) {real, imag} */,
  {32'h4270d975, 32'h41fe95b4} /* (9, 20, 8) {real, imag} */,
  {32'hc1a36cb9, 32'h42185782} /* (9, 20, 7) {real, imag} */,
  {32'h42f8b1cc, 32'h4189f9e3} /* (9, 20, 6) {real, imag} */,
  {32'h429fae32, 32'h42019336} /* (9, 20, 5) {real, imag} */,
  {32'hc3316a45, 32'h424c269c} /* (9, 20, 4) {real, imag} */,
  {32'h41862aa4, 32'hc316a083} /* (9, 20, 3) {real, imag} */,
  {32'h43fa8a88, 32'h43772e4f} /* (9, 20, 2) {real, imag} */,
  {32'hc4a37382, 32'hc2e5c240} /* (9, 20, 1) {real, imag} */,
  {32'hc40b07e4, 32'h00000000} /* (9, 20, 0) {real, imag} */,
  {32'hc5272452, 32'h433ed0e0} /* (9, 19, 31) {real, imag} */,
  {32'h448fe2b7, 32'hc3cbe218} /* (9, 19, 30) {real, imag} */,
  {32'hc2567e2a, 32'h43322659} /* (9, 19, 29) {real, imag} */,
  {32'hc3452e81, 32'h4227d064} /* (9, 19, 28) {real, imag} */,
  {32'h4304a652, 32'h41a8e4e0} /* (9, 19, 27) {real, imag} */,
  {32'h4288525e, 32'hc2d57f85} /* (9, 19, 26) {real, imag} */,
  {32'hc1b647e4, 32'h430e37cc} /* (9, 19, 25) {real, imag} */,
  {32'h42c87466, 32'hc1c7a30a} /* (9, 19, 24) {real, imag} */,
  {32'h42901333, 32'hc147d4f7} /* (9, 19, 23) {real, imag} */,
  {32'h41c9289c, 32'hc18b9112} /* (9, 19, 22) {real, imag} */,
  {32'h41898176, 32'hc2a5c2e4} /* (9, 19, 21) {real, imag} */,
  {32'hbe914c20, 32'h4245e7eb} /* (9, 19, 20) {real, imag} */,
  {32'hc27063f0, 32'h407995c0} /* (9, 19, 19) {real, imag} */,
  {32'h43020ba5, 32'hc251f142} /* (9, 19, 18) {real, imag} */,
  {32'hc0dd8d80, 32'hc09b74e9} /* (9, 19, 17) {real, imag} */,
  {32'hc10210c1, 32'h00000000} /* (9, 19, 16) {real, imag} */,
  {32'hc0dd8d80, 32'h409b74e9} /* (9, 19, 15) {real, imag} */,
  {32'h43020ba5, 32'h4251f142} /* (9, 19, 14) {real, imag} */,
  {32'hc27063f0, 32'hc07995c0} /* (9, 19, 13) {real, imag} */,
  {32'hbe914c20, 32'hc245e7eb} /* (9, 19, 12) {real, imag} */,
  {32'h41898176, 32'h42a5c2e4} /* (9, 19, 11) {real, imag} */,
  {32'h41c9289c, 32'h418b9112} /* (9, 19, 10) {real, imag} */,
  {32'h42901333, 32'h4147d4f7} /* (9, 19, 9) {real, imag} */,
  {32'h42c87466, 32'h41c7a30a} /* (9, 19, 8) {real, imag} */,
  {32'hc1b647e4, 32'hc30e37cc} /* (9, 19, 7) {real, imag} */,
  {32'h4288525e, 32'h42d57f85} /* (9, 19, 6) {real, imag} */,
  {32'h4304a652, 32'hc1a8e4e0} /* (9, 19, 5) {real, imag} */,
  {32'hc3452e81, 32'hc227d064} /* (9, 19, 4) {real, imag} */,
  {32'hc2567e2a, 32'hc3322659} /* (9, 19, 3) {real, imag} */,
  {32'h448fe2b7, 32'h43cbe218} /* (9, 19, 2) {real, imag} */,
  {32'hc5272452, 32'hc33ed0e0} /* (9, 19, 1) {real, imag} */,
  {32'hc4e0c5c5, 32'h00000000} /* (9, 19, 0) {real, imag} */,
  {32'hc566e06f, 32'h43ad142e} /* (9, 18, 31) {real, imag} */,
  {32'h44a8d5ff, 32'hc3b9d92a} /* (9, 18, 30) {real, imag} */,
  {32'hc293c72e, 32'h42aa07df} /* (9, 18, 29) {real, imag} */,
  {32'hc3762732, 32'hc1240844} /* (9, 18, 28) {real, imag} */,
  {32'h436a8c94, 32'h428ce85c} /* (9, 18, 27) {real, imag} */,
  {32'h42baeeb1, 32'hc1a18c39} /* (9, 18, 26) {real, imag} */,
  {32'hc30895f8, 32'h41b3528e} /* (9, 18, 25) {real, imag} */,
  {32'h42a77fe6, 32'hc2116aec} /* (9, 18, 24) {real, imag} */,
  {32'hc2af005e, 32'h4212cbd2} /* (9, 18, 23) {real, imag} */,
  {32'h42a5da0c, 32'h418db913} /* (9, 18, 22) {real, imag} */,
  {32'hc2999b3b, 32'hc2a458ce} /* (9, 18, 21) {real, imag} */,
  {32'h41b9fdd1, 32'h40228280} /* (9, 18, 20) {real, imag} */,
  {32'h420cbebe, 32'h415e2fd2} /* (9, 18, 19) {real, imag} */,
  {32'h420ebcfe, 32'hc241cd1c} /* (9, 18, 18) {real, imag} */,
  {32'hc116614b, 32'h421ce820} /* (9, 18, 17) {real, imag} */,
  {32'h42da3e37, 32'h00000000} /* (9, 18, 16) {real, imag} */,
  {32'hc116614b, 32'hc21ce820} /* (9, 18, 15) {real, imag} */,
  {32'h420ebcfe, 32'h4241cd1c} /* (9, 18, 14) {real, imag} */,
  {32'h420cbebe, 32'hc15e2fd2} /* (9, 18, 13) {real, imag} */,
  {32'h41b9fdd1, 32'hc0228280} /* (9, 18, 12) {real, imag} */,
  {32'hc2999b3b, 32'h42a458ce} /* (9, 18, 11) {real, imag} */,
  {32'h42a5da0c, 32'hc18db913} /* (9, 18, 10) {real, imag} */,
  {32'hc2af005e, 32'hc212cbd2} /* (9, 18, 9) {real, imag} */,
  {32'h42a77fe6, 32'h42116aec} /* (9, 18, 8) {real, imag} */,
  {32'hc30895f8, 32'hc1b3528e} /* (9, 18, 7) {real, imag} */,
  {32'h42baeeb1, 32'h41a18c39} /* (9, 18, 6) {real, imag} */,
  {32'h436a8c94, 32'hc28ce85c} /* (9, 18, 5) {real, imag} */,
  {32'hc3762732, 32'h41240844} /* (9, 18, 4) {real, imag} */,
  {32'hc293c72e, 32'hc2aa07df} /* (9, 18, 3) {real, imag} */,
  {32'h44a8d5ff, 32'h43b9d92a} /* (9, 18, 2) {real, imag} */,
  {32'hc566e06f, 32'hc3ad142e} /* (9, 18, 1) {real, imag} */,
  {32'hc51f64db, 32'h00000000} /* (9, 18, 0) {real, imag} */,
  {32'hc584309d, 32'h43b52f12} /* (9, 17, 31) {real, imag} */,
  {32'h44ba857c, 32'hc320febc} /* (9, 17, 30) {real, imag} */,
  {32'h42312796, 32'hc131789c} /* (9, 17, 29) {real, imag} */,
  {32'hc36b7fa4, 32'h41c23568} /* (9, 17, 28) {real, imag} */,
  {32'h43a03589, 32'hc17e4fc8} /* (9, 17, 27) {real, imag} */,
  {32'h4314972c, 32'hc23584fc} /* (9, 17, 26) {real, imag} */,
  {32'hc2b4fd3c, 32'hc073e148} /* (9, 17, 25) {real, imag} */,
  {32'h42a37f7a, 32'h409c7380} /* (9, 17, 24) {real, imag} */,
  {32'h42816b0a, 32'hc0ac6252} /* (9, 17, 23) {real, imag} */,
  {32'h42ea3f92, 32'h42d1bd02} /* (9, 17, 22) {real, imag} */,
  {32'hc1c31c2a, 32'hc2145b63} /* (9, 17, 21) {real, imag} */,
  {32'hc2a37095, 32'h4257b479} /* (9, 17, 20) {real, imag} */,
  {32'h427ff9d2, 32'h40f17276} /* (9, 17, 19) {real, imag} */,
  {32'hc1f9906c, 32'hc22ddc2c} /* (9, 17, 18) {real, imag} */,
  {32'h41e823e6, 32'h41178544} /* (9, 17, 17) {real, imag} */,
  {32'hc28a4bae, 32'h00000000} /* (9, 17, 16) {real, imag} */,
  {32'h41e823e6, 32'hc1178544} /* (9, 17, 15) {real, imag} */,
  {32'hc1f9906c, 32'h422ddc2c} /* (9, 17, 14) {real, imag} */,
  {32'h427ff9d2, 32'hc0f17276} /* (9, 17, 13) {real, imag} */,
  {32'hc2a37095, 32'hc257b479} /* (9, 17, 12) {real, imag} */,
  {32'hc1c31c2a, 32'h42145b63} /* (9, 17, 11) {real, imag} */,
  {32'h42ea3f92, 32'hc2d1bd02} /* (9, 17, 10) {real, imag} */,
  {32'h42816b0a, 32'h40ac6252} /* (9, 17, 9) {real, imag} */,
  {32'h42a37f7a, 32'hc09c7380} /* (9, 17, 8) {real, imag} */,
  {32'hc2b4fd3c, 32'h4073e148} /* (9, 17, 7) {real, imag} */,
  {32'h4314972c, 32'h423584fc} /* (9, 17, 6) {real, imag} */,
  {32'h43a03589, 32'h417e4fc8} /* (9, 17, 5) {real, imag} */,
  {32'hc36b7fa4, 32'hc1c23568} /* (9, 17, 4) {real, imag} */,
  {32'h42312796, 32'h4131789c} /* (9, 17, 3) {real, imag} */,
  {32'h44ba857c, 32'h4320febc} /* (9, 17, 2) {real, imag} */,
  {32'hc584309d, 32'hc3b52f12} /* (9, 17, 1) {real, imag} */,
  {32'hc54fec68, 32'h00000000} /* (9, 17, 0) {real, imag} */,
  {32'hc589f147, 32'h43b6035c} /* (9, 16, 31) {real, imag} */,
  {32'h44c68b90, 32'hc319f3d0} /* (9, 16, 30) {real, imag} */,
  {32'hc23a3a3a, 32'h41ec0622} /* (9, 16, 29) {real, imag} */,
  {32'hc295ea78, 32'h42185666} /* (9, 16, 28) {real, imag} */,
  {32'h4380b7cd, 32'hc28857f2} /* (9, 16, 27) {real, imag} */,
  {32'h43068dce, 32'hc190ca5a} /* (9, 16, 26) {real, imag} */,
  {32'hc133a02c, 32'h41f2d110} /* (9, 16, 25) {real, imag} */,
  {32'h42a4d2ec, 32'h41e32173} /* (9, 16, 24) {real, imag} */,
  {32'h42157c90, 32'h41548940} /* (9, 16, 23) {real, imag} */,
  {32'h40cd0af0, 32'hbf8fc700} /* (9, 16, 22) {real, imag} */,
  {32'h42a0df65, 32'h421d7b33} /* (9, 16, 21) {real, imag} */,
  {32'hc0a745a8, 32'hc25bb5fa} /* (9, 16, 20) {real, imag} */,
  {32'hc1eaf7ea, 32'hc2adea93} /* (9, 16, 19) {real, imag} */,
  {32'h4101b3e1, 32'hc28734ae} /* (9, 16, 18) {real, imag} */,
  {32'hc1c3a9d6, 32'hc1a1dd61} /* (9, 16, 17) {real, imag} */,
  {32'h41117098, 32'h00000000} /* (9, 16, 16) {real, imag} */,
  {32'hc1c3a9d6, 32'h41a1dd61} /* (9, 16, 15) {real, imag} */,
  {32'h4101b3e1, 32'h428734ae} /* (9, 16, 14) {real, imag} */,
  {32'hc1eaf7ea, 32'h42adea93} /* (9, 16, 13) {real, imag} */,
  {32'hc0a745a8, 32'h425bb5fa} /* (9, 16, 12) {real, imag} */,
  {32'h42a0df65, 32'hc21d7b33} /* (9, 16, 11) {real, imag} */,
  {32'h40cd0af0, 32'h3f8fc700} /* (9, 16, 10) {real, imag} */,
  {32'h42157c90, 32'hc1548940} /* (9, 16, 9) {real, imag} */,
  {32'h42a4d2ec, 32'hc1e32173} /* (9, 16, 8) {real, imag} */,
  {32'hc133a02c, 32'hc1f2d110} /* (9, 16, 7) {real, imag} */,
  {32'h43068dce, 32'h4190ca5a} /* (9, 16, 6) {real, imag} */,
  {32'h4380b7cd, 32'h428857f2} /* (9, 16, 5) {real, imag} */,
  {32'hc295ea78, 32'hc2185666} /* (9, 16, 4) {real, imag} */,
  {32'hc23a3a3a, 32'hc1ec0622} /* (9, 16, 3) {real, imag} */,
  {32'h44c68b90, 32'h4319f3d0} /* (9, 16, 2) {real, imag} */,
  {32'hc589f147, 32'hc3b6035c} /* (9, 16, 1) {real, imag} */,
  {32'hc557fb42, 32'h00000000} /* (9, 16, 0) {real, imag} */,
  {32'hc5894b6b, 32'h43a2746e} /* (9, 15, 31) {real, imag} */,
  {32'h44c30904, 32'hc351fb8c} /* (9, 15, 30) {real, imag} */,
  {32'h40eaa870, 32'hc14476dc} /* (9, 15, 29) {real, imag} */,
  {32'hc35d7316, 32'h4212ee20} /* (9, 15, 28) {real, imag} */,
  {32'h4329d75a, 32'hc2e9a025} /* (9, 15, 27) {real, imag} */,
  {32'h42badbdf, 32'h41c72a1f} /* (9, 15, 26) {real, imag} */,
  {32'hc201ec4c, 32'hc10ff8a6} /* (9, 15, 25) {real, imag} */,
  {32'h42d1c740, 32'h41a3ba88} /* (9, 15, 24) {real, imag} */,
  {32'hc1f367ef, 32'h416e3deb} /* (9, 15, 23) {real, imag} */,
  {32'hc09e77f8, 32'hc25583b0} /* (9, 15, 22) {real, imag} */,
  {32'h41c90d3c, 32'hc1bc3204} /* (9, 15, 21) {real, imag} */,
  {32'hc228822e, 32'hc27f6437} /* (9, 15, 20) {real, imag} */,
  {32'hc2731b4e, 32'hc08a9446} /* (9, 15, 19) {real, imag} */,
  {32'h412e5f21, 32'hc10b017c} /* (9, 15, 18) {real, imag} */,
  {32'hc22d4c11, 32'h4222ede9} /* (9, 15, 17) {real, imag} */,
  {32'hc23886f0, 32'h00000000} /* (9, 15, 16) {real, imag} */,
  {32'hc22d4c11, 32'hc222ede9} /* (9, 15, 15) {real, imag} */,
  {32'h412e5f21, 32'h410b017c} /* (9, 15, 14) {real, imag} */,
  {32'hc2731b4e, 32'h408a9446} /* (9, 15, 13) {real, imag} */,
  {32'hc228822e, 32'h427f6437} /* (9, 15, 12) {real, imag} */,
  {32'h41c90d3c, 32'h41bc3204} /* (9, 15, 11) {real, imag} */,
  {32'hc09e77f8, 32'h425583b0} /* (9, 15, 10) {real, imag} */,
  {32'hc1f367ef, 32'hc16e3deb} /* (9, 15, 9) {real, imag} */,
  {32'h42d1c740, 32'hc1a3ba88} /* (9, 15, 8) {real, imag} */,
  {32'hc201ec4c, 32'h410ff8a6} /* (9, 15, 7) {real, imag} */,
  {32'h42badbdf, 32'hc1c72a1f} /* (9, 15, 6) {real, imag} */,
  {32'h4329d75a, 32'h42e9a025} /* (9, 15, 5) {real, imag} */,
  {32'hc35d7316, 32'hc212ee20} /* (9, 15, 4) {real, imag} */,
  {32'h40eaa870, 32'h414476dc} /* (9, 15, 3) {real, imag} */,
  {32'h44c30904, 32'h4351fb8c} /* (9, 15, 2) {real, imag} */,
  {32'hc5894b6b, 32'hc3a2746e} /* (9, 15, 1) {real, imag} */,
  {32'hc54f7f1e, 32'h00000000} /* (9, 15, 0) {real, imag} */,
  {32'hc57884bb, 32'h43ba7cba} /* (9, 14, 31) {real, imag} */,
  {32'h44b70375, 32'hc34445cc} /* (9, 14, 30) {real, imag} */,
  {32'h42cafb5a, 32'h4305e0ce} /* (9, 14, 29) {real, imag} */,
  {32'hc38ada2d, 32'hc2958b78} /* (9, 14, 28) {real, imag} */,
  {32'h431a1c74, 32'hc2fe884e} /* (9, 14, 27) {real, imag} */,
  {32'hc1e173d8, 32'h4255c078} /* (9, 14, 26) {real, imag} */,
  {32'hc1bf42fc, 32'h42587d97} /* (9, 14, 25) {real, imag} */,
  {32'h42e626f4, 32'h422dbfd4} /* (9, 14, 24) {real, imag} */,
  {32'h42a57774, 32'hc2552b1e} /* (9, 14, 23) {real, imag} */,
  {32'h42eea30e, 32'h4259d7fe} /* (9, 14, 22) {real, imag} */,
  {32'h4255ea3a, 32'hc289da0a} /* (9, 14, 21) {real, imag} */,
  {32'hc033a5c8, 32'hc28fc69c} /* (9, 14, 20) {real, imag} */,
  {32'hc210a58e, 32'h419b266b} /* (9, 14, 19) {real, imag} */,
  {32'hc223ff82, 32'h40e7c3f0} /* (9, 14, 18) {real, imag} */,
  {32'h410a5101, 32'h4273c104} /* (9, 14, 17) {real, imag} */,
  {32'h429a0625, 32'h00000000} /* (9, 14, 16) {real, imag} */,
  {32'h410a5101, 32'hc273c104} /* (9, 14, 15) {real, imag} */,
  {32'hc223ff82, 32'hc0e7c3f0} /* (9, 14, 14) {real, imag} */,
  {32'hc210a58e, 32'hc19b266b} /* (9, 14, 13) {real, imag} */,
  {32'hc033a5c8, 32'h428fc69c} /* (9, 14, 12) {real, imag} */,
  {32'h4255ea3a, 32'h4289da0a} /* (9, 14, 11) {real, imag} */,
  {32'h42eea30e, 32'hc259d7fe} /* (9, 14, 10) {real, imag} */,
  {32'h42a57774, 32'h42552b1e} /* (9, 14, 9) {real, imag} */,
  {32'h42e626f4, 32'hc22dbfd4} /* (9, 14, 8) {real, imag} */,
  {32'hc1bf42fc, 32'hc2587d97} /* (9, 14, 7) {real, imag} */,
  {32'hc1e173d8, 32'hc255c078} /* (9, 14, 6) {real, imag} */,
  {32'h431a1c74, 32'h42fe884e} /* (9, 14, 5) {real, imag} */,
  {32'hc38ada2d, 32'h42958b78} /* (9, 14, 4) {real, imag} */,
  {32'h42cafb5a, 32'hc305e0ce} /* (9, 14, 3) {real, imag} */,
  {32'h44b70375, 32'h434445cc} /* (9, 14, 2) {real, imag} */,
  {32'hc57884bb, 32'hc3ba7cba} /* (9, 14, 1) {real, imag} */,
  {32'hc53d213d, 32'h00000000} /* (9, 14, 0) {real, imag} */,
  {32'hc550853c, 32'h4269cf40} /* (9, 13, 31) {real, imag} */,
  {32'h449f7c6f, 32'hc307e30f} /* (9, 13, 30) {real, imag} */,
  {32'h424d6604, 32'h4299b7a4} /* (9, 13, 29) {real, imag} */,
  {32'hc39b4d73, 32'h41aed904} /* (9, 13, 28) {real, imag} */,
  {32'h4369bf32, 32'hc2d9af50} /* (9, 13, 27) {real, imag} */,
  {32'h41330bec, 32'h423e8036} /* (9, 13, 26) {real, imag} */,
  {32'hc286f44f, 32'hc1cd7898} /* (9, 13, 25) {real, imag} */,
  {32'hc206940b, 32'h416d6244} /* (9, 13, 24) {real, imag} */,
  {32'hc26da4a6, 32'hc202a95f} /* (9, 13, 23) {real, imag} */,
  {32'hc2c0fbf9, 32'h41feb312} /* (9, 13, 22) {real, imag} */,
  {32'h4122650b, 32'hc197f8df} /* (9, 13, 21) {real, imag} */,
  {32'h41d03ffe, 32'hc12b8dc0} /* (9, 13, 20) {real, imag} */,
  {32'h410d3d02, 32'h427d2d06} /* (9, 13, 19) {real, imag} */,
  {32'hc249ac04, 32'hc3277fbe} /* (9, 13, 18) {real, imag} */,
  {32'hc08e8c58, 32'hc1877abc} /* (9, 13, 17) {real, imag} */,
  {32'h4202d54c, 32'h00000000} /* (9, 13, 16) {real, imag} */,
  {32'hc08e8c58, 32'h41877abc} /* (9, 13, 15) {real, imag} */,
  {32'hc249ac04, 32'h43277fbe} /* (9, 13, 14) {real, imag} */,
  {32'h410d3d02, 32'hc27d2d06} /* (9, 13, 13) {real, imag} */,
  {32'h41d03ffe, 32'h412b8dc0} /* (9, 13, 12) {real, imag} */,
  {32'h4122650b, 32'h4197f8df} /* (9, 13, 11) {real, imag} */,
  {32'hc2c0fbf9, 32'hc1feb312} /* (9, 13, 10) {real, imag} */,
  {32'hc26da4a6, 32'h4202a95f} /* (9, 13, 9) {real, imag} */,
  {32'hc206940b, 32'hc16d6244} /* (9, 13, 8) {real, imag} */,
  {32'hc286f44f, 32'h41cd7898} /* (9, 13, 7) {real, imag} */,
  {32'h41330bec, 32'hc23e8036} /* (9, 13, 6) {real, imag} */,
  {32'h4369bf32, 32'h42d9af50} /* (9, 13, 5) {real, imag} */,
  {32'hc39b4d73, 32'hc1aed904} /* (9, 13, 4) {real, imag} */,
  {32'h424d6604, 32'hc299b7a4} /* (9, 13, 3) {real, imag} */,
  {32'h449f7c6f, 32'h4307e30f} /* (9, 13, 2) {real, imag} */,
  {32'hc550853c, 32'hc269cf40} /* (9, 13, 1) {real, imag} */,
  {32'hc51d934e, 32'h00000000} /* (9, 13, 0) {real, imag} */,
  {32'hc51b21bd, 32'hc3182a20} /* (9, 12, 31) {real, imag} */,
  {32'h44802ff8, 32'h3fc5e980} /* (9, 12, 30) {real, imag} */,
  {32'h425cfbc8, 32'h42af0064} /* (9, 12, 29) {real, imag} */,
  {32'hc33a18f3, 32'h419018b8} /* (9, 12, 28) {real, imag} */,
  {32'h431ba2fd, 32'hc0d548bc} /* (9, 12, 27) {real, imag} */,
  {32'h41b68cbe, 32'hc0d720eb} /* (9, 12, 26) {real, imag} */,
  {32'hc28ac006, 32'h41164af8} /* (9, 12, 25) {real, imag} */,
  {32'h42ea11b2, 32'hc274ba7c} /* (9, 12, 24) {real, imag} */,
  {32'hc0c936f8, 32'h42866a7e} /* (9, 12, 23) {real, imag} */,
  {32'hc253f10c, 32'h407a2860} /* (9, 12, 22) {real, imag} */,
  {32'hc1af45f5, 32'hc2c247c2} /* (9, 12, 21) {real, imag} */,
  {32'h4161e4b3, 32'hc15a961f} /* (9, 12, 20) {real, imag} */,
  {32'hc15d1a08, 32'hc21859c4} /* (9, 12, 19) {real, imag} */,
  {32'hc13d7185, 32'h429bd703} /* (9, 12, 18) {real, imag} */,
  {32'hc2474adc, 32'hc28c1302} /* (9, 12, 17) {real, imag} */,
  {32'h41468bc0, 32'h00000000} /* (9, 12, 16) {real, imag} */,
  {32'hc2474adc, 32'h428c1302} /* (9, 12, 15) {real, imag} */,
  {32'hc13d7185, 32'hc29bd703} /* (9, 12, 14) {real, imag} */,
  {32'hc15d1a08, 32'h421859c4} /* (9, 12, 13) {real, imag} */,
  {32'h4161e4b3, 32'h415a961f} /* (9, 12, 12) {real, imag} */,
  {32'hc1af45f5, 32'h42c247c2} /* (9, 12, 11) {real, imag} */,
  {32'hc253f10c, 32'hc07a2860} /* (9, 12, 10) {real, imag} */,
  {32'hc0c936f8, 32'hc2866a7e} /* (9, 12, 9) {real, imag} */,
  {32'h42ea11b2, 32'h4274ba7c} /* (9, 12, 8) {real, imag} */,
  {32'hc28ac006, 32'hc1164af8} /* (9, 12, 7) {real, imag} */,
  {32'h41b68cbe, 32'h40d720eb} /* (9, 12, 6) {real, imag} */,
  {32'h431ba2fd, 32'h40d548bc} /* (9, 12, 5) {real, imag} */,
  {32'hc33a18f3, 32'hc19018b8} /* (9, 12, 4) {real, imag} */,
  {32'h425cfbc8, 32'hc2af0064} /* (9, 12, 3) {real, imag} */,
  {32'h44802ff8, 32'hbfc5e980} /* (9, 12, 2) {real, imag} */,
  {32'hc51b21bd, 32'h43182a20} /* (9, 12, 1) {real, imag} */,
  {32'hc4d33986, 32'h00000000} /* (9, 12, 0) {real, imag} */,
  {32'hc48c5114, 32'hc3938701} /* (9, 11, 31) {real, imag} */,
  {32'h44099b16, 32'h423b8b44} /* (9, 11, 30) {real, imag} */,
  {32'hbfb67c10, 32'h41b40ec4} /* (9, 11, 29) {real, imag} */,
  {32'hc3011512, 32'hc30f88f6} /* (9, 11, 28) {real, imag} */,
  {32'h428c9572, 32'hc18f8462} /* (9, 11, 27) {real, imag} */,
  {32'hc193d1ae, 32'hc2b1cc2c} /* (9, 11, 26) {real, imag} */,
  {32'h41f5768c, 32'hc21f2b26} /* (9, 11, 25) {real, imag} */,
  {32'h42481aca, 32'h414f6468} /* (9, 11, 24) {real, imag} */,
  {32'hc224a900, 32'hbf361ee0} /* (9, 11, 23) {real, imag} */,
  {32'h42bbea08, 32'hc24de2d7} /* (9, 11, 22) {real, imag} */,
  {32'h429478b3, 32'hc2f45568} /* (9, 11, 21) {real, imag} */,
  {32'hc21363ae, 32'h41854b68} /* (9, 11, 20) {real, imag} */,
  {32'h41a9120f, 32'h3f6fa5c0} /* (9, 11, 19) {real, imag} */,
  {32'h41be9340, 32'h41d07624} /* (9, 11, 18) {real, imag} */,
  {32'hc1497cc1, 32'h4243a168} /* (9, 11, 17) {real, imag} */,
  {32'h4262814f, 32'h00000000} /* (9, 11, 16) {real, imag} */,
  {32'hc1497cc1, 32'hc243a168} /* (9, 11, 15) {real, imag} */,
  {32'h41be9340, 32'hc1d07624} /* (9, 11, 14) {real, imag} */,
  {32'h41a9120f, 32'hbf6fa5c0} /* (9, 11, 13) {real, imag} */,
  {32'hc21363ae, 32'hc1854b68} /* (9, 11, 12) {real, imag} */,
  {32'h429478b3, 32'h42f45568} /* (9, 11, 11) {real, imag} */,
  {32'h42bbea08, 32'h424de2d7} /* (9, 11, 10) {real, imag} */,
  {32'hc224a900, 32'h3f361ee0} /* (9, 11, 9) {real, imag} */,
  {32'h42481aca, 32'hc14f6468} /* (9, 11, 8) {real, imag} */,
  {32'h41f5768c, 32'h421f2b26} /* (9, 11, 7) {real, imag} */,
  {32'hc193d1ae, 32'h42b1cc2c} /* (9, 11, 6) {real, imag} */,
  {32'h428c9572, 32'h418f8462} /* (9, 11, 5) {real, imag} */,
  {32'hc3011512, 32'h430f88f6} /* (9, 11, 4) {real, imag} */,
  {32'hbfb67c10, 32'hc1b40ec4} /* (9, 11, 3) {real, imag} */,
  {32'h44099b16, 32'hc23b8b44} /* (9, 11, 2) {real, imag} */,
  {32'hc48c5114, 32'h43938701} /* (9, 11, 1) {real, imag} */,
  {32'hc3b98164, 32'h00000000} /* (9, 11, 0) {real, imag} */,
  {32'h442794d0, 32'hc431adf4} /* (9, 10, 31) {real, imag} */,
  {32'hc38c58d0, 32'h43631598} /* (9, 10, 30) {real, imag} */,
  {32'hc22a1340, 32'hc232bdca} /* (9, 10, 29) {real, imag} */,
  {32'hc2a5390d, 32'hc37ff851} /* (9, 10, 28) {real, imag} */,
  {32'hc2be68b2, 32'h3f2a2060} /* (9, 10, 27) {real, imag} */,
  {32'h42f69ab2, 32'h41589b60} /* (9, 10, 26) {real, imag} */,
  {32'h4230f37a, 32'hc1b3c6d0} /* (9, 10, 25) {real, imag} */,
  {32'hc0e36392, 32'h428a400e} /* (9, 10, 24) {real, imag} */,
  {32'h41f53065, 32'hbff15780} /* (9, 10, 23) {real, imag} */,
  {32'h428e4de1, 32'h3ee48240} /* (9, 10, 22) {real, imag} */,
  {32'hc0c98cf8, 32'hc24604ff} /* (9, 10, 21) {real, imag} */,
  {32'h41a76d8e, 32'h425d0ec4} /* (9, 10, 20) {real, imag} */,
  {32'h42d8d4d0, 32'hc2ac1d36} /* (9, 10, 19) {real, imag} */,
  {32'hc249184c, 32'hc2917e4e} /* (9, 10, 18) {real, imag} */,
  {32'h4203582c, 32'h4223d38a} /* (9, 10, 17) {real, imag} */,
  {32'hc2f6bf91, 32'h00000000} /* (9, 10, 16) {real, imag} */,
  {32'h4203582c, 32'hc223d38a} /* (9, 10, 15) {real, imag} */,
  {32'hc249184c, 32'h42917e4e} /* (9, 10, 14) {real, imag} */,
  {32'h42d8d4d0, 32'h42ac1d36} /* (9, 10, 13) {real, imag} */,
  {32'h41a76d8e, 32'hc25d0ec4} /* (9, 10, 12) {real, imag} */,
  {32'hc0c98cf8, 32'h424604ff} /* (9, 10, 11) {real, imag} */,
  {32'h428e4de1, 32'hbee48240} /* (9, 10, 10) {real, imag} */,
  {32'h41f53065, 32'h3ff15780} /* (9, 10, 9) {real, imag} */,
  {32'hc0e36392, 32'hc28a400e} /* (9, 10, 8) {real, imag} */,
  {32'h4230f37a, 32'h41b3c6d0} /* (9, 10, 7) {real, imag} */,
  {32'h42f69ab2, 32'hc1589b60} /* (9, 10, 6) {real, imag} */,
  {32'hc2be68b2, 32'hbf2a2060} /* (9, 10, 5) {real, imag} */,
  {32'hc2a5390d, 32'h437ff851} /* (9, 10, 4) {real, imag} */,
  {32'hc22a1340, 32'h4232bdca} /* (9, 10, 3) {real, imag} */,
  {32'hc38c58d0, 32'hc3631598} /* (9, 10, 2) {real, imag} */,
  {32'h442794d0, 32'h4431adf4} /* (9, 10, 1) {real, imag} */,
  {32'h449007bf, 32'h00000000} /* (9, 10, 0) {real, imag} */,
  {32'h45004fee, 32'hc496357a} /* (9, 9, 31) {real, imag} */,
  {32'hc447ceac, 32'h43c96ce2} /* (9, 9, 30) {real, imag} */,
  {32'hc232fc59, 32'hc22f1dae} /* (9, 9, 29) {real, imag} */,
  {32'hc2863fa9, 32'hc347883e} /* (9, 9, 28) {real, imag} */,
  {32'hc323305e, 32'h429f57bc} /* (9, 9, 27) {real, imag} */,
  {32'h423ef7d0, 32'hc246bb24} /* (9, 9, 26) {real, imag} */,
  {32'h412983c8, 32'h42d4505c} /* (9, 9, 25) {real, imag} */,
  {32'hc18075e5, 32'hc1b3343a} /* (9, 9, 24) {real, imag} */,
  {32'hc24a1383, 32'hc246254d} /* (9, 9, 23) {real, imag} */,
  {32'hc0c9b016, 32'h417ae2a6} /* (9, 9, 22) {real, imag} */,
  {32'hc1496098, 32'h3f097940} /* (9, 9, 21) {real, imag} */,
  {32'h428e516a, 32'h409b5580} /* (9, 9, 20) {real, imag} */,
  {32'h41829270, 32'hc13498e4} /* (9, 9, 19) {real, imag} */,
  {32'h4177a500, 32'h424f69bc} /* (9, 9, 18) {real, imag} */,
  {32'h404cdef0, 32'hc20dc564} /* (9, 9, 17) {real, imag} */,
  {32'hc2765732, 32'h00000000} /* (9, 9, 16) {real, imag} */,
  {32'h404cdef0, 32'h420dc564} /* (9, 9, 15) {real, imag} */,
  {32'h4177a500, 32'hc24f69bc} /* (9, 9, 14) {real, imag} */,
  {32'h41829270, 32'h413498e4} /* (9, 9, 13) {real, imag} */,
  {32'h428e516a, 32'hc09b5580} /* (9, 9, 12) {real, imag} */,
  {32'hc1496098, 32'hbf097940} /* (9, 9, 11) {real, imag} */,
  {32'hc0c9b016, 32'hc17ae2a6} /* (9, 9, 10) {real, imag} */,
  {32'hc24a1383, 32'h4246254d} /* (9, 9, 9) {real, imag} */,
  {32'hc18075e5, 32'h41b3343a} /* (9, 9, 8) {real, imag} */,
  {32'h412983c8, 32'hc2d4505c} /* (9, 9, 7) {real, imag} */,
  {32'h423ef7d0, 32'h4246bb24} /* (9, 9, 6) {real, imag} */,
  {32'hc323305e, 32'hc29f57bc} /* (9, 9, 5) {real, imag} */,
  {32'hc2863fa9, 32'h4347883e} /* (9, 9, 4) {real, imag} */,
  {32'hc232fc59, 32'h422f1dae} /* (9, 9, 3) {real, imag} */,
  {32'hc447ceac, 32'hc3c96ce2} /* (9, 9, 2) {real, imag} */,
  {32'h45004fee, 32'h4496357a} /* (9, 9, 1) {real, imag} */,
  {32'h450f9792, 32'h00000000} /* (9, 9, 0) {real, imag} */,
  {32'h4534b00a, 32'hc4b8b947} /* (9, 8, 31) {real, imag} */,
  {32'hc48f078d, 32'h440d2a50} /* (9, 8, 30) {real, imag} */,
  {32'hc290f7b8, 32'hc2fb2505} /* (9, 8, 29) {real, imag} */,
  {32'h4218ed98, 32'hc32143fd} /* (9, 8, 28) {real, imag} */,
  {32'hc2fc382a, 32'h4299327d} /* (9, 8, 27) {real, imag} */,
  {32'hc287426d, 32'h429de48b} /* (9, 8, 26) {real, imag} */,
  {32'h42413866, 32'h4226dda8} /* (9, 8, 25) {real, imag} */,
  {32'hc25bdf2c, 32'hc24866bc} /* (9, 8, 24) {real, imag} */,
  {32'h41655bbe, 32'h4118d644} /* (9, 8, 23) {real, imag} */,
  {32'h422c7e88, 32'h41ebeed4} /* (9, 8, 22) {real, imag} */,
  {32'hc2421fcc, 32'h42037388} /* (9, 8, 21) {real, imag} */,
  {32'h41969688, 32'hc1bdefac} /* (9, 8, 20) {real, imag} */,
  {32'hc1d44678, 32'hc276fd0a} /* (9, 8, 19) {real, imag} */,
  {32'hc26a4a1e, 32'hc1878b84} /* (9, 8, 18) {real, imag} */,
  {32'hc1ac05dc, 32'hc2894762} /* (9, 8, 17) {real, imag} */,
  {32'hc20725b6, 32'h00000000} /* (9, 8, 16) {real, imag} */,
  {32'hc1ac05dc, 32'h42894762} /* (9, 8, 15) {real, imag} */,
  {32'hc26a4a1e, 32'h41878b84} /* (9, 8, 14) {real, imag} */,
  {32'hc1d44678, 32'h4276fd0a} /* (9, 8, 13) {real, imag} */,
  {32'h41969688, 32'h41bdefac} /* (9, 8, 12) {real, imag} */,
  {32'hc2421fcc, 32'hc2037388} /* (9, 8, 11) {real, imag} */,
  {32'h422c7e88, 32'hc1ebeed4} /* (9, 8, 10) {real, imag} */,
  {32'h41655bbe, 32'hc118d644} /* (9, 8, 9) {real, imag} */,
  {32'hc25bdf2c, 32'h424866bc} /* (9, 8, 8) {real, imag} */,
  {32'h42413866, 32'hc226dda8} /* (9, 8, 7) {real, imag} */,
  {32'hc287426d, 32'hc29de48b} /* (9, 8, 6) {real, imag} */,
  {32'hc2fc382a, 32'hc299327d} /* (9, 8, 5) {real, imag} */,
  {32'h4218ed98, 32'h432143fd} /* (9, 8, 4) {real, imag} */,
  {32'hc290f7b8, 32'h42fb2505} /* (9, 8, 3) {real, imag} */,
  {32'hc48f078d, 32'hc40d2a50} /* (9, 8, 2) {real, imag} */,
  {32'h4534b00a, 32'h44b8b947} /* (9, 8, 1) {real, imag} */,
  {32'h455a19f1, 32'h00000000} /* (9, 8, 0) {real, imag} */,
  {32'h45564cfd, 32'hc4e449ee} /* (9, 7, 31) {real, imag} */,
  {32'hc48c9735, 32'h444da56b} /* (9, 7, 30) {real, imag} */,
  {32'hc20349c9, 32'hc2d57579} /* (9, 7, 29) {real, imag} */,
  {32'h42c55541, 32'hc28d00ae} /* (9, 7, 28) {real, imag} */,
  {32'hc35e3930, 32'h43436732} /* (9, 7, 27) {real, imag} */,
  {32'hbca7c000, 32'h413f0a09} /* (9, 7, 26) {real, imag} */,
  {32'h42ca47b2, 32'h420af8d0} /* (9, 7, 25) {real, imag} */,
  {32'hc1819245, 32'h426d5eed} /* (9, 7, 24) {real, imag} */,
  {32'h41ad86a3, 32'h4276d93c} /* (9, 7, 23) {real, imag} */,
  {32'h4263bac5, 32'h3f46c780} /* (9, 7, 22) {real, imag} */,
  {32'hc2689952, 32'h41ca84cf} /* (9, 7, 21) {real, imag} */,
  {32'hc20c6e9e, 32'hc23e1232} /* (9, 7, 20) {real, imag} */,
  {32'hc289f0eb, 32'hc1b2549a} /* (9, 7, 19) {real, imag} */,
  {32'h421cb390, 32'hc2266042} /* (9, 7, 18) {real, imag} */,
  {32'hc0943d26, 32'h419bb0cd} /* (9, 7, 17) {real, imag} */,
  {32'h425fa17a, 32'h00000000} /* (9, 7, 16) {real, imag} */,
  {32'hc0943d26, 32'hc19bb0cd} /* (9, 7, 15) {real, imag} */,
  {32'h421cb390, 32'h42266042} /* (9, 7, 14) {real, imag} */,
  {32'hc289f0eb, 32'h41b2549a} /* (9, 7, 13) {real, imag} */,
  {32'hc20c6e9e, 32'h423e1232} /* (9, 7, 12) {real, imag} */,
  {32'hc2689952, 32'hc1ca84cf} /* (9, 7, 11) {real, imag} */,
  {32'h4263bac5, 32'hbf46c780} /* (9, 7, 10) {real, imag} */,
  {32'h41ad86a3, 32'hc276d93c} /* (9, 7, 9) {real, imag} */,
  {32'hc1819245, 32'hc26d5eed} /* (9, 7, 8) {real, imag} */,
  {32'h42ca47b2, 32'hc20af8d0} /* (9, 7, 7) {real, imag} */,
  {32'hbca7c000, 32'hc13f0a09} /* (9, 7, 6) {real, imag} */,
  {32'hc35e3930, 32'hc3436732} /* (9, 7, 5) {real, imag} */,
  {32'h42c55541, 32'h428d00ae} /* (9, 7, 4) {real, imag} */,
  {32'hc20349c9, 32'h42d57579} /* (9, 7, 3) {real, imag} */,
  {32'hc48c9735, 32'hc44da56b} /* (9, 7, 2) {real, imag} */,
  {32'h45564cfd, 32'h44e449ee} /* (9, 7, 1) {real, imag} */,
  {32'h45845442, 32'h00000000} /* (9, 7, 0) {real, imag} */,
  {32'h4562b082, 32'hc5150e2e} /* (9, 6, 31) {real, imag} */,
  {32'hc46c602d, 32'h4484e77d} /* (9, 6, 30) {real, imag} */,
  {32'hc1c81b89, 32'hc1474bd0} /* (9, 6, 29) {real, imag} */,
  {32'h423b0b1e, 32'hc2b2d53e} /* (9, 6, 28) {real, imag} */,
  {32'hc33a53f2, 32'h423518b2} /* (9, 6, 27) {real, imag} */,
  {32'h425b1e4c, 32'h42ae7a2d} /* (9, 6, 26) {real, imag} */,
  {32'h4306bac6, 32'h42f7ca74} /* (9, 6, 25) {real, imag} */,
  {32'h41f1715c, 32'h42b5601f} /* (9, 6, 24) {real, imag} */,
  {32'hc21de3ba, 32'hc12152f1} /* (9, 6, 23) {real, imag} */,
  {32'hc19a3c35, 32'h423758a0} /* (9, 6, 22) {real, imag} */,
  {32'h3cacf000, 32'hc26b3009} /* (9, 6, 21) {real, imag} */,
  {32'h4000a1d4, 32'hc231df62} /* (9, 6, 20) {real, imag} */,
  {32'h41aad3da, 32'hc24f4764} /* (9, 6, 19) {real, imag} */,
  {32'h4252dc52, 32'h42d403d9} /* (9, 6, 18) {real, imag} */,
  {32'hc27aa253, 32'h42193a38} /* (9, 6, 17) {real, imag} */,
  {32'hc2baeaf4, 32'h00000000} /* (9, 6, 16) {real, imag} */,
  {32'hc27aa253, 32'hc2193a38} /* (9, 6, 15) {real, imag} */,
  {32'h4252dc52, 32'hc2d403d9} /* (9, 6, 14) {real, imag} */,
  {32'h41aad3da, 32'h424f4764} /* (9, 6, 13) {real, imag} */,
  {32'h4000a1d4, 32'h4231df62} /* (9, 6, 12) {real, imag} */,
  {32'h3cacf000, 32'h426b3009} /* (9, 6, 11) {real, imag} */,
  {32'hc19a3c35, 32'hc23758a0} /* (9, 6, 10) {real, imag} */,
  {32'hc21de3ba, 32'h412152f1} /* (9, 6, 9) {real, imag} */,
  {32'h41f1715c, 32'hc2b5601f} /* (9, 6, 8) {real, imag} */,
  {32'h4306bac6, 32'hc2f7ca74} /* (9, 6, 7) {real, imag} */,
  {32'h425b1e4c, 32'hc2ae7a2d} /* (9, 6, 6) {real, imag} */,
  {32'hc33a53f2, 32'hc23518b2} /* (9, 6, 5) {real, imag} */,
  {32'h423b0b1e, 32'h42b2d53e} /* (9, 6, 4) {real, imag} */,
  {32'hc1c81b89, 32'h41474bd0} /* (9, 6, 3) {real, imag} */,
  {32'hc46c602d, 32'hc484e77d} /* (9, 6, 2) {real, imag} */,
  {32'h4562b082, 32'h45150e2e} /* (9, 6, 1) {real, imag} */,
  {32'h45960f59, 32'h00000000} /* (9, 6, 0) {real, imag} */,
  {32'h455ab55d, 32'hc5423622} /* (9, 5, 31) {real, imag} */,
  {32'hc3bf16b0, 32'h449f2cf6} /* (9, 5, 30) {real, imag} */,
  {32'hc2c725ab, 32'h419f7c46} /* (9, 5, 29) {real, imag} */,
  {32'h4101e020, 32'h42335bf8} /* (9, 5, 28) {real, imag} */,
  {32'hc26e26eb, 32'h42a3ed8d} /* (9, 5, 27) {real, imag} */,
  {32'h42fb3226, 32'h42ad268c} /* (9, 5, 26) {real, imag} */,
  {32'h4255bf41, 32'hc05a6bc0} /* (9, 5, 25) {real, imag} */,
  {32'hc1e4cbb7, 32'h4300563b} /* (9, 5, 24) {real, imag} */,
  {32'hc2ad3a05, 32'hc2c4d508} /* (9, 5, 23) {real, imag} */,
  {32'h42ec3cf2, 32'h42801e58} /* (9, 5, 22) {real, imag} */,
  {32'h42854d29, 32'hc2ccf716} /* (9, 5, 21) {real, imag} */,
  {32'hc12dd86a, 32'h414ce108} /* (9, 5, 20) {real, imag} */,
  {32'h423e7e1d, 32'h42ce61c2} /* (9, 5, 19) {real, imag} */,
  {32'hc2c5acf6, 32'h42ef20f2} /* (9, 5, 18) {real, imag} */,
  {32'h4115b5dc, 32'h41fb4ea1} /* (9, 5, 17) {real, imag} */,
  {32'h4202c51d, 32'h00000000} /* (9, 5, 16) {real, imag} */,
  {32'h4115b5dc, 32'hc1fb4ea1} /* (9, 5, 15) {real, imag} */,
  {32'hc2c5acf6, 32'hc2ef20f2} /* (9, 5, 14) {real, imag} */,
  {32'h423e7e1d, 32'hc2ce61c2} /* (9, 5, 13) {real, imag} */,
  {32'hc12dd86a, 32'hc14ce108} /* (9, 5, 12) {real, imag} */,
  {32'h42854d29, 32'h42ccf716} /* (9, 5, 11) {real, imag} */,
  {32'h42ec3cf2, 32'hc2801e58} /* (9, 5, 10) {real, imag} */,
  {32'hc2ad3a05, 32'h42c4d508} /* (9, 5, 9) {real, imag} */,
  {32'hc1e4cbb7, 32'hc300563b} /* (9, 5, 8) {real, imag} */,
  {32'h4255bf41, 32'h405a6bc0} /* (9, 5, 7) {real, imag} */,
  {32'h42fb3226, 32'hc2ad268c} /* (9, 5, 6) {real, imag} */,
  {32'hc26e26eb, 32'hc2a3ed8d} /* (9, 5, 5) {real, imag} */,
  {32'h4101e020, 32'hc2335bf8} /* (9, 5, 4) {real, imag} */,
  {32'hc2c725ab, 32'hc19f7c46} /* (9, 5, 3) {real, imag} */,
  {32'hc3bf16b0, 32'hc49f2cf6} /* (9, 5, 2) {real, imag} */,
  {32'h455ab55d, 32'h45423622} /* (9, 5, 1) {real, imag} */,
  {32'h45a93d4c, 32'h00000000} /* (9, 5, 0) {real, imag} */,
  {32'h4555c031, 32'hc56785f7} /* (9, 4, 31) {real, imag} */,
  {32'hc1684300, 32'h4494cf60} /* (9, 4, 30) {real, imag} */,
  {32'hc2b3a628, 32'hc22d1e07} /* (9, 4, 29) {real, imag} */,
  {32'hc27ff010, 32'h437bf1c4} /* (9, 4, 28) {real, imag} */,
  {32'hc2f82f00, 32'h42f981fd} /* (9, 4, 27) {real, imag} */,
  {32'hc15eadf4, 32'hc29595c4} /* (9, 4, 26) {real, imag} */,
  {32'h4317f305, 32'hc2bac1f6} /* (9, 4, 25) {real, imag} */,
  {32'hc0810372, 32'hc093cdea} /* (9, 4, 24) {real, imag} */,
  {32'hc1e8ba76, 32'hc1649b28} /* (9, 4, 23) {real, imag} */,
  {32'h41c6f99a, 32'h43095548} /* (9, 4, 22) {real, imag} */,
  {32'hc2318527, 32'hc23be2c9} /* (9, 4, 21) {real, imag} */,
  {32'h421aab88, 32'hc13fc873} /* (9, 4, 20) {real, imag} */,
  {32'h4270faa8, 32'hc2a6643a} /* (9, 4, 19) {real, imag} */,
  {32'h419009ce, 32'hc297856e} /* (9, 4, 18) {real, imag} */,
  {32'hc1a660e6, 32'h42374277} /* (9, 4, 17) {real, imag} */,
  {32'hc193fedc, 32'h00000000} /* (9, 4, 16) {real, imag} */,
  {32'hc1a660e6, 32'hc2374277} /* (9, 4, 15) {real, imag} */,
  {32'h419009ce, 32'h4297856e} /* (9, 4, 14) {real, imag} */,
  {32'h4270faa8, 32'h42a6643a} /* (9, 4, 13) {real, imag} */,
  {32'h421aab88, 32'h413fc873} /* (9, 4, 12) {real, imag} */,
  {32'hc2318527, 32'h423be2c9} /* (9, 4, 11) {real, imag} */,
  {32'h41c6f99a, 32'hc3095548} /* (9, 4, 10) {real, imag} */,
  {32'hc1e8ba76, 32'h41649b28} /* (9, 4, 9) {real, imag} */,
  {32'hc0810372, 32'h4093cdea} /* (9, 4, 8) {real, imag} */,
  {32'h4317f305, 32'h42bac1f6} /* (9, 4, 7) {real, imag} */,
  {32'hc15eadf4, 32'h429595c4} /* (9, 4, 6) {real, imag} */,
  {32'hc2f82f00, 32'hc2f981fd} /* (9, 4, 5) {real, imag} */,
  {32'hc27ff010, 32'hc37bf1c4} /* (9, 4, 4) {real, imag} */,
  {32'hc2b3a628, 32'h422d1e07} /* (9, 4, 3) {real, imag} */,
  {32'hc1684300, 32'hc494cf60} /* (9, 4, 2) {real, imag} */,
  {32'h4555c031, 32'h456785f7} /* (9, 4, 1) {real, imag} */,
  {32'h45b017fc, 32'h00000000} /* (9, 4, 0) {real, imag} */,
  {32'h454f4f16, 32'hc57c4646} /* (9, 3, 31) {real, imag} */,
  {32'h439fdaac, 32'h4494d3fe} /* (9, 3, 30) {real, imag} */,
  {32'hc2dd6987, 32'h42e0ea11} /* (9, 3, 29) {real, imag} */,
  {32'hc2831a84, 32'h438b0ab6} /* (9, 3, 28) {real, imag} */,
  {32'hc2c47331, 32'h41ff5061} /* (9, 3, 27) {real, imag} */,
  {32'hc25414f7, 32'hc280938a} /* (9, 3, 26) {real, imag} */,
  {32'h42da9a8f, 32'h41963374} /* (9, 3, 25) {real, imag} */,
  {32'h415211ab, 32'h4335bb5c} /* (9, 3, 24) {real, imag} */,
  {32'hc25f4b0b, 32'h4175f3aa} /* (9, 3, 23) {real, imag} */,
  {32'h42666fc2, 32'h42d24c2a} /* (9, 3, 22) {real, imag} */,
  {32'hc0ac11c8, 32'h4280fec6} /* (9, 3, 21) {real, imag} */,
  {32'h42287f36, 32'h41fa3cf4} /* (9, 3, 20) {real, imag} */,
  {32'h41ed4479, 32'h42814574} /* (9, 3, 19) {real, imag} */,
  {32'h41cf821b, 32'h41ef474f} /* (9, 3, 18) {real, imag} */,
  {32'hc2946d96, 32'hc22dd8f0} /* (9, 3, 17) {real, imag} */,
  {32'h41f2f514, 32'h00000000} /* (9, 3, 16) {real, imag} */,
  {32'hc2946d96, 32'h422dd8f0} /* (9, 3, 15) {real, imag} */,
  {32'h41cf821b, 32'hc1ef474f} /* (9, 3, 14) {real, imag} */,
  {32'h41ed4479, 32'hc2814574} /* (9, 3, 13) {real, imag} */,
  {32'h42287f36, 32'hc1fa3cf4} /* (9, 3, 12) {real, imag} */,
  {32'hc0ac11c8, 32'hc280fec6} /* (9, 3, 11) {real, imag} */,
  {32'h42666fc2, 32'hc2d24c2a} /* (9, 3, 10) {real, imag} */,
  {32'hc25f4b0b, 32'hc175f3aa} /* (9, 3, 9) {real, imag} */,
  {32'h415211ab, 32'hc335bb5c} /* (9, 3, 8) {real, imag} */,
  {32'h42da9a8f, 32'hc1963374} /* (9, 3, 7) {real, imag} */,
  {32'hc25414f7, 32'h4280938a} /* (9, 3, 6) {real, imag} */,
  {32'hc2c47331, 32'hc1ff5061} /* (9, 3, 5) {real, imag} */,
  {32'hc2831a84, 32'hc38b0ab6} /* (9, 3, 4) {real, imag} */,
  {32'hc2dd6987, 32'hc2e0ea11} /* (9, 3, 3) {real, imag} */,
  {32'h439fdaac, 32'hc494d3fe} /* (9, 3, 2) {real, imag} */,
  {32'h454f4f16, 32'h457c4646} /* (9, 3, 1) {real, imag} */,
  {32'h45b2f865, 32'h00000000} /* (9, 3, 0) {real, imag} */,
  {32'h45440347, 32'hc57b92e6} /* (9, 2, 31) {real, imag} */,
  {32'h43b803f1, 32'h44893b88} /* (9, 2, 30) {real, imag} */,
  {32'hc35e44bc, 32'h432aa7a6} /* (9, 2, 29) {real, imag} */,
  {32'hc19cb78c, 32'h43971dd4} /* (9, 2, 28) {real, imag} */,
  {32'hc2b9fc36, 32'hc356e856} /* (9, 2, 27) {real, imag} */,
  {32'hc2f845ae, 32'hc21959d0} /* (9, 2, 26) {real, imag} */,
  {32'h4136eeaa, 32'hc1897cc6} /* (9, 2, 25) {real, imag} */,
  {32'h42a746d9, 32'h42e9171a} /* (9, 2, 24) {real, imag} */,
  {32'hc118ce58, 32'h4015f2b2} /* (9, 2, 23) {real, imag} */,
  {32'hc2e0d2d1, 32'h423f2510} /* (9, 2, 22) {real, imag} */,
  {32'hc2ecaffe, 32'hc2b67f2a} /* (9, 2, 21) {real, imag} */,
  {32'h423885f4, 32'h42379a7a} /* (9, 2, 20) {real, imag} */,
  {32'h423d7be2, 32'hc2ac1ade} /* (9, 2, 19) {real, imag} */,
  {32'hc16a9578, 32'h41f84ce4} /* (9, 2, 18) {real, imag} */,
  {32'hc0996587, 32'h41e05a3a} /* (9, 2, 17) {real, imag} */,
  {32'h4220d688, 32'h00000000} /* (9, 2, 16) {real, imag} */,
  {32'hc0996587, 32'hc1e05a3a} /* (9, 2, 15) {real, imag} */,
  {32'hc16a9578, 32'hc1f84ce4} /* (9, 2, 14) {real, imag} */,
  {32'h423d7be2, 32'h42ac1ade} /* (9, 2, 13) {real, imag} */,
  {32'h423885f4, 32'hc2379a7a} /* (9, 2, 12) {real, imag} */,
  {32'hc2ecaffe, 32'h42b67f2a} /* (9, 2, 11) {real, imag} */,
  {32'hc2e0d2d1, 32'hc23f2510} /* (9, 2, 10) {real, imag} */,
  {32'hc118ce58, 32'hc015f2b2} /* (9, 2, 9) {real, imag} */,
  {32'h42a746d9, 32'hc2e9171a} /* (9, 2, 8) {real, imag} */,
  {32'h4136eeaa, 32'h41897cc6} /* (9, 2, 7) {real, imag} */,
  {32'hc2f845ae, 32'h421959d0} /* (9, 2, 6) {real, imag} */,
  {32'hc2b9fc36, 32'h4356e856} /* (9, 2, 5) {real, imag} */,
  {32'hc19cb78c, 32'hc3971dd4} /* (9, 2, 4) {real, imag} */,
  {32'hc35e44bc, 32'hc32aa7a6} /* (9, 2, 3) {real, imag} */,
  {32'h43b803f1, 32'hc4893b88} /* (9, 2, 2) {real, imag} */,
  {32'h45440347, 32'h457b92e6} /* (9, 2, 1) {real, imag} */,
  {32'h45b61095, 32'h00000000} /* (9, 2, 0) {real, imag} */,
  {32'h454fb855, 32'hc56a1c71} /* (9, 1, 31) {real, imag} */,
  {32'h4387ba5c, 32'h447f7470} /* (9, 1, 30) {real, imag} */,
  {32'hc39f3bc5, 32'h422be16b} /* (9, 1, 29) {real, imag} */,
  {32'h40f1e3c8, 32'h43a60387} /* (9, 1, 28) {real, imag} */,
  {32'hc3234561, 32'hc3303336} /* (9, 1, 27) {real, imag} */,
  {32'hc1efc840, 32'h421ed080} /* (9, 1, 26) {real, imag} */,
  {32'h414d7d12, 32'h4173f18a} /* (9, 1, 25) {real, imag} */,
  {32'h427f6b28, 32'h42897cae} /* (9, 1, 24) {real, imag} */,
  {32'h42333654, 32'hc1caba62} /* (9, 1, 23) {real, imag} */,
  {32'hc29b90f2, 32'hbfb9dba8} /* (9, 1, 22) {real, imag} */,
  {32'hc291280c, 32'hbf8b0100} /* (9, 1, 21) {real, imag} */,
  {32'h419c0964, 32'h42a4a1b2} /* (9, 1, 20) {real, imag} */,
  {32'h42c1a4ae, 32'hc2b80ef8} /* (9, 1, 19) {real, imag} */,
  {32'hc2017487, 32'h41c1a182} /* (9, 1, 18) {real, imag} */,
  {32'hc0c71a93, 32'hc20693f4} /* (9, 1, 17) {real, imag} */,
  {32'hc1d820bf, 32'h00000000} /* (9, 1, 16) {real, imag} */,
  {32'hc0c71a93, 32'h420693f4} /* (9, 1, 15) {real, imag} */,
  {32'hc2017487, 32'hc1c1a182} /* (9, 1, 14) {real, imag} */,
  {32'h42c1a4ae, 32'h42b80ef8} /* (9, 1, 13) {real, imag} */,
  {32'h419c0964, 32'hc2a4a1b2} /* (9, 1, 12) {real, imag} */,
  {32'hc291280c, 32'h3f8b0100} /* (9, 1, 11) {real, imag} */,
  {32'hc29b90f2, 32'h3fb9dba8} /* (9, 1, 10) {real, imag} */,
  {32'h42333654, 32'h41caba62} /* (9, 1, 9) {real, imag} */,
  {32'h427f6b28, 32'hc2897cae} /* (9, 1, 8) {real, imag} */,
  {32'h414d7d12, 32'hc173f18a} /* (9, 1, 7) {real, imag} */,
  {32'hc1efc840, 32'hc21ed080} /* (9, 1, 6) {real, imag} */,
  {32'hc3234561, 32'h43303336} /* (9, 1, 5) {real, imag} */,
  {32'h40f1e3c8, 32'hc3a60387} /* (9, 1, 4) {real, imag} */,
  {32'hc39f3bc5, 32'hc22be16b} /* (9, 1, 3) {real, imag} */,
  {32'h4387ba5c, 32'hc47f7470} /* (9, 1, 2) {real, imag} */,
  {32'h454fb855, 32'h456a1c71} /* (9, 1, 1) {real, imag} */,
  {32'h45b359c9, 32'h00000000} /* (9, 1, 0) {real, imag} */,
  {32'h455d1b56, 32'hc53c6bd6} /* (9, 0, 31) {real, imag} */,
  {32'hc3163e04, 32'h4457a754} /* (9, 0, 30) {real, imag} */,
  {32'hc343f42c, 32'h4282e6e4} /* (9, 0, 29) {real, imag} */,
  {32'h42623904, 32'h43134cf0} /* (9, 0, 28) {real, imag} */,
  {32'hc2de8181, 32'hc2b3078c} /* (9, 0, 27) {real, imag} */,
  {32'h41e772b8, 32'hc1edf8c6} /* (9, 0, 26) {real, imag} */,
  {32'h41b94da8, 32'h40856962} /* (9, 0, 25) {real, imag} */,
  {32'hbf664840, 32'hc1df6d81} /* (9, 0, 24) {real, imag} */,
  {32'h411bf2e4, 32'hc23ad7d2} /* (9, 0, 23) {real, imag} */,
  {32'hc2597e8b, 32'hc107d0e0} /* (9, 0, 22) {real, imag} */,
  {32'hc1c73cb8, 32'h4234c8f7} /* (9, 0, 21) {real, imag} */,
  {32'hc20a114d, 32'h41c4ea0f} /* (9, 0, 20) {real, imag} */,
  {32'hc23ba99d, 32'h4235328a} /* (9, 0, 19) {real, imag} */,
  {32'h416ee83d, 32'h41e5c313} /* (9, 0, 18) {real, imag} */,
  {32'hc1b105f2, 32'hc1ded6a3} /* (9, 0, 17) {real, imag} */,
  {32'h42993aa9, 32'h00000000} /* (9, 0, 16) {real, imag} */,
  {32'hc1b105f2, 32'h41ded6a3} /* (9, 0, 15) {real, imag} */,
  {32'h416ee83d, 32'hc1e5c313} /* (9, 0, 14) {real, imag} */,
  {32'hc23ba99d, 32'hc235328a} /* (9, 0, 13) {real, imag} */,
  {32'hc20a114d, 32'hc1c4ea0f} /* (9, 0, 12) {real, imag} */,
  {32'hc1c73cb8, 32'hc234c8f7} /* (9, 0, 11) {real, imag} */,
  {32'hc2597e8b, 32'h4107d0e0} /* (9, 0, 10) {real, imag} */,
  {32'h411bf2e4, 32'h423ad7d2} /* (9, 0, 9) {real, imag} */,
  {32'hbf664840, 32'h41df6d81} /* (9, 0, 8) {real, imag} */,
  {32'h41b94da8, 32'hc0856962} /* (9, 0, 7) {real, imag} */,
  {32'h41e772b8, 32'h41edf8c6} /* (9, 0, 6) {real, imag} */,
  {32'hc2de8181, 32'h42b3078c} /* (9, 0, 5) {real, imag} */,
  {32'h42623904, 32'hc3134cf0} /* (9, 0, 4) {real, imag} */,
  {32'hc343f42c, 32'hc282e6e4} /* (9, 0, 3) {real, imag} */,
  {32'hc3163e04, 32'hc457a754} /* (9, 0, 2) {real, imag} */,
  {32'h455d1b56, 32'h453c6bd6} /* (9, 0, 1) {real, imag} */,
  {32'h45a8b349, 32'h00000000} /* (9, 0, 0) {real, imag} */,
  {32'h4562e33d, 32'hc4fb271c} /* (8, 31, 31) {real, imag} */,
  {32'hc43667ba, 32'h440b375e} /* (8, 31, 30) {real, imag} */,
  {32'hc237a3d2, 32'hc1fb6b58} /* (8, 31, 29) {real, imag} */,
  {32'h41b90f2e, 32'h42c57365} /* (8, 31, 28) {real, imag} */,
  {32'hc303a102, 32'h4045dea0} /* (8, 31, 27) {real, imag} */,
  {32'h40e687ec, 32'hbe8a67c0} /* (8, 31, 26) {real, imag} */,
  {32'h427baa56, 32'hbee9c680} /* (8, 31, 25) {real, imag} */,
  {32'hc2c699a0, 32'h41b8d2eb} /* (8, 31, 24) {real, imag} */,
  {32'h4294bc9e, 32'hc15de536} /* (8, 31, 23) {real, imag} */,
  {32'h42ba5c88, 32'h415acaa4} /* (8, 31, 22) {real, imag} */,
  {32'hc25094f3, 32'h428f8234} /* (8, 31, 21) {real, imag} */,
  {32'hc238766b, 32'hc23ae02e} /* (8, 31, 20) {real, imag} */,
  {32'h42581694, 32'hc209cc5c} /* (8, 31, 19) {real, imag} */,
  {32'hc22ac209, 32'h4210e7d9} /* (8, 31, 18) {real, imag} */,
  {32'hc1e21969, 32'hc281f6d5} /* (8, 31, 17) {real, imag} */,
  {32'h423e4c6f, 32'h00000000} /* (8, 31, 16) {real, imag} */,
  {32'hc1e21969, 32'h4281f6d5} /* (8, 31, 15) {real, imag} */,
  {32'hc22ac209, 32'hc210e7d9} /* (8, 31, 14) {real, imag} */,
  {32'h42581694, 32'h4209cc5c} /* (8, 31, 13) {real, imag} */,
  {32'hc238766b, 32'h423ae02e} /* (8, 31, 12) {real, imag} */,
  {32'hc25094f3, 32'hc28f8234} /* (8, 31, 11) {real, imag} */,
  {32'h42ba5c88, 32'hc15acaa4} /* (8, 31, 10) {real, imag} */,
  {32'h4294bc9e, 32'h415de536} /* (8, 31, 9) {real, imag} */,
  {32'hc2c699a0, 32'hc1b8d2eb} /* (8, 31, 8) {real, imag} */,
  {32'h427baa56, 32'h3ee9c680} /* (8, 31, 7) {real, imag} */,
  {32'h40e687ec, 32'h3e8a67c0} /* (8, 31, 6) {real, imag} */,
  {32'hc303a102, 32'hc045dea0} /* (8, 31, 5) {real, imag} */,
  {32'h41b90f2e, 32'hc2c57365} /* (8, 31, 4) {real, imag} */,
  {32'hc237a3d2, 32'h41fb6b58} /* (8, 31, 3) {real, imag} */,
  {32'hc43667ba, 32'hc40b375e} /* (8, 31, 2) {real, imag} */,
  {32'h4562e33d, 32'h44fb271c} /* (8, 31, 1) {real, imag} */,
  {32'h45a28aaf, 32'h00000000} /* (8, 31, 0) {real, imag} */,
  {32'h4582e612, 32'hc4c58433} /* (8, 30, 31) {real, imag} */,
  {32'hc488f4f1, 32'h4403e919} /* (8, 30, 30) {real, imag} */,
  {32'h3fa73080, 32'h422c57f6} /* (8, 30, 29) {real, imag} */,
  {32'h42491036, 32'h407c5680} /* (8, 30, 28) {real, imag} */,
  {32'hc32a107a, 32'h42994a9a} /* (8, 30, 27) {real, imag} */,
  {32'h42d608e8, 32'h41c813c5} /* (8, 30, 26) {real, imag} */,
  {32'h429ddf37, 32'hc185a42e} /* (8, 30, 25) {real, imag} */,
  {32'hc2b81ea0, 32'h43242dfc} /* (8, 30, 24) {real, imag} */,
  {32'h429090aa, 32'hc1ded204} /* (8, 30, 23) {real, imag} */,
  {32'hc303626a, 32'h40348a00} /* (8, 30, 22) {real, imag} */,
  {32'hc31da687, 32'h4250b30c} /* (8, 30, 21) {real, imag} */,
  {32'hc25266d0, 32'hc14a75cc} /* (8, 30, 20) {real, imag} */,
  {32'h42aa3318, 32'h40e15f00} /* (8, 30, 19) {real, imag} */,
  {32'hc26ae84e, 32'h429db482} /* (8, 30, 18) {real, imag} */,
  {32'hc20ac3c9, 32'hc0679340} /* (8, 30, 17) {real, imag} */,
  {32'hc1a8afa8, 32'h00000000} /* (8, 30, 16) {real, imag} */,
  {32'hc20ac3c9, 32'h40679340} /* (8, 30, 15) {real, imag} */,
  {32'hc26ae84e, 32'hc29db482} /* (8, 30, 14) {real, imag} */,
  {32'h42aa3318, 32'hc0e15f00} /* (8, 30, 13) {real, imag} */,
  {32'hc25266d0, 32'h414a75cc} /* (8, 30, 12) {real, imag} */,
  {32'hc31da687, 32'hc250b30c} /* (8, 30, 11) {real, imag} */,
  {32'hc303626a, 32'hc0348a00} /* (8, 30, 10) {real, imag} */,
  {32'h429090aa, 32'h41ded204} /* (8, 30, 9) {real, imag} */,
  {32'hc2b81ea0, 32'hc3242dfc} /* (8, 30, 8) {real, imag} */,
  {32'h429ddf37, 32'h4185a42e} /* (8, 30, 7) {real, imag} */,
  {32'h42d608e8, 32'hc1c813c5} /* (8, 30, 6) {real, imag} */,
  {32'hc32a107a, 32'hc2994a9a} /* (8, 30, 5) {real, imag} */,
  {32'h42491036, 32'hc07c5680} /* (8, 30, 4) {real, imag} */,
  {32'h3fa73080, 32'hc22c57f6} /* (8, 30, 3) {real, imag} */,
  {32'hc488f4f1, 32'hc403e919} /* (8, 30, 2) {real, imag} */,
  {32'h4582e612, 32'h44c58433} /* (8, 30, 1) {real, imag} */,
  {32'h45a839b4, 32'h00000000} /* (8, 30, 0) {real, imag} */,
  {32'h458d906c, 32'hc493c068} /* (8, 29, 31) {real, imag} */,
  {32'hc49012aa, 32'h44028db4} /* (8, 29, 30) {real, imag} */,
  {32'h42cf5cd2, 32'h42a3ab9c} /* (8, 29, 29) {real, imag} */,
  {32'h43472fce, 32'hc2685edc} /* (8, 29, 28) {real, imag} */,
  {32'hc37033c6, 32'h42a73851} /* (8, 29, 27) {real, imag} */,
  {32'h41ca5b3c, 32'hbf3e5e00} /* (8, 29, 26) {real, imag} */,
  {32'h419b9c30, 32'hc2b569d1} /* (8, 29, 25) {real, imag} */,
  {32'hc2e2d9fb, 32'h429d1f3a} /* (8, 29, 24) {real, imag} */,
  {32'hc217088d, 32'h41f0026a} /* (8, 29, 23) {real, imag} */,
  {32'hc25beb76, 32'hc1984a82} /* (8, 29, 22) {real, imag} */,
  {32'hc3060289, 32'h424113ee} /* (8, 29, 21) {real, imag} */,
  {32'hc089e7a0, 32'h41327023} /* (8, 29, 20) {real, imag} */,
  {32'hc0cf79f0, 32'hc21410b1} /* (8, 29, 19) {real, imag} */,
  {32'hc1f45e70, 32'h42e0a1de} /* (8, 29, 18) {real, imag} */,
  {32'hc1710870, 32'hc20a2d3d} /* (8, 29, 17) {real, imag} */,
  {32'hc19444a8, 32'h00000000} /* (8, 29, 16) {real, imag} */,
  {32'hc1710870, 32'h420a2d3d} /* (8, 29, 15) {real, imag} */,
  {32'hc1f45e70, 32'hc2e0a1de} /* (8, 29, 14) {real, imag} */,
  {32'hc0cf79f0, 32'h421410b1} /* (8, 29, 13) {real, imag} */,
  {32'hc089e7a0, 32'hc1327023} /* (8, 29, 12) {real, imag} */,
  {32'hc3060289, 32'hc24113ee} /* (8, 29, 11) {real, imag} */,
  {32'hc25beb76, 32'h41984a82} /* (8, 29, 10) {real, imag} */,
  {32'hc217088d, 32'hc1f0026a} /* (8, 29, 9) {real, imag} */,
  {32'hc2e2d9fb, 32'hc29d1f3a} /* (8, 29, 8) {real, imag} */,
  {32'h419b9c30, 32'h42b569d1} /* (8, 29, 7) {real, imag} */,
  {32'h41ca5b3c, 32'h3f3e5e00} /* (8, 29, 6) {real, imag} */,
  {32'hc37033c6, 32'hc2a73851} /* (8, 29, 5) {real, imag} */,
  {32'h43472fce, 32'h42685edc} /* (8, 29, 4) {real, imag} */,
  {32'h42cf5cd2, 32'hc2a3ab9c} /* (8, 29, 3) {real, imag} */,
  {32'hc49012aa, 32'hc4028db4} /* (8, 29, 2) {real, imag} */,
  {32'h458d906c, 32'h4493c068} /* (8, 29, 1) {real, imag} */,
  {32'h45a1f8d5, 32'h00000000} /* (8, 29, 0) {real, imag} */,
  {32'h458f57ae, 32'hc47a587e} /* (8, 28, 31) {real, imag} */,
  {32'hc4abf274, 32'h44149a39} /* (8, 28, 30) {real, imag} */,
  {32'h40d99c80, 32'hc09f6960} /* (8, 28, 29) {real, imag} */,
  {32'h435bad6c, 32'hbe5af000} /* (8, 28, 28) {real, imag} */,
  {32'hc3687df2, 32'h4109b428} /* (8, 28, 27) {real, imag} */,
  {32'hc244a29c, 32'hc2696e54} /* (8, 28, 26) {real, imag} */,
  {32'hc290b664, 32'hc306073f} /* (8, 28, 25) {real, imag} */,
  {32'hc250ddb6, 32'h42a89302} /* (8, 28, 24) {real, imag} */,
  {32'hc29db5a2, 32'h4296d644} /* (8, 28, 23) {real, imag} */,
  {32'hc1f8e43e, 32'hc1eed1f8} /* (8, 28, 22) {real, imag} */,
  {32'h4160ad34, 32'h415dc080} /* (8, 28, 21) {real, imag} */,
  {32'hc22565c7, 32'hc1f0b88c} /* (8, 28, 20) {real, imag} */,
  {32'h423775fa, 32'h3f41baa0} /* (8, 28, 19) {real, imag} */,
  {32'hc20b8600, 32'h41d401d4} /* (8, 28, 18) {real, imag} */,
  {32'h42d1f7fe, 32'hc2f95b36} /* (8, 28, 17) {real, imag} */,
  {32'h427f3cb4, 32'h00000000} /* (8, 28, 16) {real, imag} */,
  {32'h42d1f7fe, 32'h42f95b36} /* (8, 28, 15) {real, imag} */,
  {32'hc20b8600, 32'hc1d401d4} /* (8, 28, 14) {real, imag} */,
  {32'h423775fa, 32'hbf41baa0} /* (8, 28, 13) {real, imag} */,
  {32'hc22565c7, 32'h41f0b88c} /* (8, 28, 12) {real, imag} */,
  {32'h4160ad34, 32'hc15dc080} /* (8, 28, 11) {real, imag} */,
  {32'hc1f8e43e, 32'h41eed1f8} /* (8, 28, 10) {real, imag} */,
  {32'hc29db5a2, 32'hc296d644} /* (8, 28, 9) {real, imag} */,
  {32'hc250ddb6, 32'hc2a89302} /* (8, 28, 8) {real, imag} */,
  {32'hc290b664, 32'h4306073f} /* (8, 28, 7) {real, imag} */,
  {32'hc244a29c, 32'h42696e54} /* (8, 28, 6) {real, imag} */,
  {32'hc3687df2, 32'hc109b428} /* (8, 28, 5) {real, imag} */,
  {32'h435bad6c, 32'h3e5af000} /* (8, 28, 4) {real, imag} */,
  {32'h40d99c80, 32'h409f6960} /* (8, 28, 3) {real, imag} */,
  {32'hc4abf274, 32'hc4149a39} /* (8, 28, 2) {real, imag} */,
  {32'h458f57ae, 32'h447a587e} /* (8, 28, 1) {real, imag} */,
  {32'h459dec2e, 32'h00000000} /* (8, 28, 0) {real, imag} */,
  {32'h45926426, 32'hc443dd94} /* (8, 27, 31) {real, imag} */,
  {32'hc4cb6a58, 32'h43ef2ebd} /* (8, 27, 30) {real, imag} */,
  {32'h42dab9de, 32'h3f9ec760} /* (8, 27, 29) {real, imag} */,
  {32'h4321aeb5, 32'hc244ce2a} /* (8, 27, 28) {real, imag} */,
  {32'hc31aa9e8, 32'h41c18861} /* (8, 27, 27) {real, imag} */,
  {32'hc228affa, 32'hc2e193d8} /* (8, 27, 26) {real, imag} */,
  {32'h42bac754, 32'hc2a941cc} /* (8, 27, 25) {real, imag} */,
  {32'h42c181d6, 32'h41a34e02} /* (8, 27, 24) {real, imag} */,
  {32'h4150b5b1, 32'h425f1546} /* (8, 27, 23) {real, imag} */,
  {32'hc02c4d20, 32'h42d0277e} /* (8, 27, 22) {real, imag} */,
  {32'hbfce3380, 32'h427e1b1c} /* (8, 27, 21) {real, imag} */,
  {32'hc2d56215, 32'hc2e34ea8} /* (8, 27, 20) {real, imag} */,
  {32'hc2efafc3, 32'h42745136} /* (8, 27, 19) {real, imag} */,
  {32'h42ad3704, 32'h41d9d4c4} /* (8, 27, 18) {real, imag} */,
  {32'h426cd9a8, 32'h412d8d80} /* (8, 27, 17) {real, imag} */,
  {32'h420f557c, 32'h00000000} /* (8, 27, 16) {real, imag} */,
  {32'h426cd9a8, 32'hc12d8d80} /* (8, 27, 15) {real, imag} */,
  {32'h42ad3704, 32'hc1d9d4c4} /* (8, 27, 14) {real, imag} */,
  {32'hc2efafc3, 32'hc2745136} /* (8, 27, 13) {real, imag} */,
  {32'hc2d56215, 32'h42e34ea8} /* (8, 27, 12) {real, imag} */,
  {32'hbfce3380, 32'hc27e1b1c} /* (8, 27, 11) {real, imag} */,
  {32'hc02c4d20, 32'hc2d0277e} /* (8, 27, 10) {real, imag} */,
  {32'h4150b5b1, 32'hc25f1546} /* (8, 27, 9) {real, imag} */,
  {32'h42c181d6, 32'hc1a34e02} /* (8, 27, 8) {real, imag} */,
  {32'h42bac754, 32'h42a941cc} /* (8, 27, 7) {real, imag} */,
  {32'hc228affa, 32'h42e193d8} /* (8, 27, 6) {real, imag} */,
  {32'hc31aa9e8, 32'hc1c18861} /* (8, 27, 5) {real, imag} */,
  {32'h4321aeb5, 32'h4244ce2a} /* (8, 27, 4) {real, imag} */,
  {32'h42dab9de, 32'hbf9ec760} /* (8, 27, 3) {real, imag} */,
  {32'hc4cb6a58, 32'hc3ef2ebd} /* (8, 27, 2) {real, imag} */,
  {32'h45926426, 32'h4443dd94} /* (8, 27, 1) {real, imag} */,
  {32'h459f0b34, 32'h00000000} /* (8, 27, 0) {real, imag} */,
  {32'h458e900d, 32'hc4133d16} /* (8, 26, 31) {real, imag} */,
  {32'hc4ce6715, 32'h439d6402} /* (8, 26, 30) {real, imag} */,
  {32'h3fc35770, 32'hc1e862d7} /* (8, 26, 29) {real, imag} */,
  {32'h437108c8, 32'h41b71eee} /* (8, 26, 28) {real, imag} */,
  {32'hc32a3011, 32'h42466871} /* (8, 26, 27) {real, imag} */,
  {32'hc2369201, 32'hc1fea270} /* (8, 26, 26) {real, imag} */,
  {32'h41b06d1c, 32'hc2e2e991} /* (8, 26, 25) {real, imag} */,
  {32'h427d9324, 32'h423341e9} /* (8, 26, 24) {real, imag} */,
  {32'h41322cc9, 32'h42a9e579} /* (8, 26, 23) {real, imag} */,
  {32'h4244881e, 32'hc1930950} /* (8, 26, 22) {real, imag} */,
  {32'hc29293ae, 32'h4159b358} /* (8, 26, 21) {real, imag} */,
  {32'hc320668e, 32'hc28ea0d0} /* (8, 26, 20) {real, imag} */,
  {32'hc2172654, 32'hc20cb08a} /* (8, 26, 19) {real, imag} */,
  {32'hc0ecf8f2, 32'h41a6966e} /* (8, 26, 18) {real, imag} */,
  {32'hc0f59810, 32'hc22f8614} /* (8, 26, 17) {real, imag} */,
  {32'h42128d78, 32'h00000000} /* (8, 26, 16) {real, imag} */,
  {32'hc0f59810, 32'h422f8614} /* (8, 26, 15) {real, imag} */,
  {32'hc0ecf8f2, 32'hc1a6966e} /* (8, 26, 14) {real, imag} */,
  {32'hc2172654, 32'h420cb08a} /* (8, 26, 13) {real, imag} */,
  {32'hc320668e, 32'h428ea0d0} /* (8, 26, 12) {real, imag} */,
  {32'hc29293ae, 32'hc159b358} /* (8, 26, 11) {real, imag} */,
  {32'h4244881e, 32'h41930950} /* (8, 26, 10) {real, imag} */,
  {32'h41322cc9, 32'hc2a9e579} /* (8, 26, 9) {real, imag} */,
  {32'h427d9324, 32'hc23341e9} /* (8, 26, 8) {real, imag} */,
  {32'h41b06d1c, 32'h42e2e991} /* (8, 26, 7) {real, imag} */,
  {32'hc2369201, 32'h41fea270} /* (8, 26, 6) {real, imag} */,
  {32'hc32a3011, 32'hc2466871} /* (8, 26, 5) {real, imag} */,
  {32'h437108c8, 32'hc1b71eee} /* (8, 26, 4) {real, imag} */,
  {32'h3fc35770, 32'h41e862d7} /* (8, 26, 3) {real, imag} */,
  {32'hc4ce6715, 32'hc39d6402} /* (8, 26, 2) {real, imag} */,
  {32'h458e900d, 32'h44133d16} /* (8, 26, 1) {real, imag} */,
  {32'h45963245, 32'h00000000} /* (8, 26, 0) {real, imag} */,
  {32'h4583c709, 32'hc3ef5d8c} /* (8, 25, 31) {real, imag} */,
  {32'hc4bc878c, 32'h4375822e} /* (8, 25, 30) {real, imag} */,
  {32'hc27d9ad1, 32'hc28f8c47} /* (8, 25, 29) {real, imag} */,
  {32'h43564962, 32'hc0a6bcd0} /* (8, 25, 28) {real, imag} */,
  {32'hc3699dc4, 32'hc1057c30} /* (8, 25, 27) {real, imag} */,
  {32'h422fa309, 32'h41bff562} /* (8, 25, 26) {real, imag} */,
  {32'hc16ab85c, 32'hc2b8861e} /* (8, 25, 25) {real, imag} */,
  {32'h4299ab00, 32'h4290883c} /* (8, 25, 24) {real, imag} */,
  {32'h41ba017c, 32'h42635a5a} /* (8, 25, 23) {real, imag} */,
  {32'hc17ad758, 32'h40e05556} /* (8, 25, 22) {real, imag} */,
  {32'hc2823736, 32'h42969b11} /* (8, 25, 21) {real, imag} */,
  {32'hc2900dea, 32'hc0fe9368} /* (8, 25, 20) {real, imag} */,
  {32'h423de1aa, 32'hc1b44361} /* (8, 25, 19) {real, imag} */,
  {32'h426397f8, 32'h41ef4196} /* (8, 25, 18) {real, imag} */,
  {32'h3f133840, 32'h416c3efa} /* (8, 25, 17) {real, imag} */,
  {32'hc1151663, 32'h00000000} /* (8, 25, 16) {real, imag} */,
  {32'h3f133840, 32'hc16c3efa} /* (8, 25, 15) {real, imag} */,
  {32'h426397f8, 32'hc1ef4196} /* (8, 25, 14) {real, imag} */,
  {32'h423de1aa, 32'h41b44361} /* (8, 25, 13) {real, imag} */,
  {32'hc2900dea, 32'h40fe9368} /* (8, 25, 12) {real, imag} */,
  {32'hc2823736, 32'hc2969b11} /* (8, 25, 11) {real, imag} */,
  {32'hc17ad758, 32'hc0e05556} /* (8, 25, 10) {real, imag} */,
  {32'h41ba017c, 32'hc2635a5a} /* (8, 25, 9) {real, imag} */,
  {32'h4299ab00, 32'hc290883c} /* (8, 25, 8) {real, imag} */,
  {32'hc16ab85c, 32'h42b8861e} /* (8, 25, 7) {real, imag} */,
  {32'h422fa309, 32'hc1bff562} /* (8, 25, 6) {real, imag} */,
  {32'hc3699dc4, 32'h41057c30} /* (8, 25, 5) {real, imag} */,
  {32'h43564962, 32'h40a6bcd0} /* (8, 25, 4) {real, imag} */,
  {32'hc27d9ad1, 32'h428f8c47} /* (8, 25, 3) {real, imag} */,
  {32'hc4bc878c, 32'hc375822e} /* (8, 25, 2) {real, imag} */,
  {32'h4583c709, 32'h43ef5d8c} /* (8, 25, 1) {real, imag} */,
  {32'h45897753, 32'h00000000} /* (8, 25, 0) {real, imag} */,
  {32'h456d9426, 32'hc3c3ce30} /* (8, 24, 31) {real, imag} */,
  {32'hc4b7431a, 32'h4322aa0a} /* (8, 24, 30) {real, imag} */,
  {32'hc2c3779d, 32'hc291a886} /* (8, 24, 29) {real, imag} */,
  {32'h43101ed8, 32'h42861a28} /* (8, 24, 28) {real, imag} */,
  {32'hc362aa3a, 32'h42df470a} /* (8, 24, 27) {real, imag} */,
  {32'h4320199c, 32'h41e4be22} /* (8, 24, 26) {real, imag} */,
  {32'hc1d5d98a, 32'hc28445f8} /* (8, 24, 25) {real, imag} */,
  {32'hc212654b, 32'h42cdb43e} /* (8, 24, 24) {real, imag} */,
  {32'h41df0b14, 32'hc2c3e2ff} /* (8, 24, 23) {real, imag} */,
  {32'h40e21b00, 32'h421ac8b2} /* (8, 24, 22) {real, imag} */,
  {32'hc29c8a2b, 32'h42236375} /* (8, 24, 21) {real, imag} */,
  {32'hc2a91fba, 32'h4293f1ff} /* (8, 24, 20) {real, imag} */,
  {32'hc2b0074c, 32'h42787344} /* (8, 24, 19) {real, imag} */,
  {32'hc0eb1ba0, 32'h416e0586} /* (8, 24, 18) {real, imag} */,
  {32'hc26c0b18, 32'h424eaed7} /* (8, 24, 17) {real, imag} */,
  {32'h42f380fb, 32'h00000000} /* (8, 24, 16) {real, imag} */,
  {32'hc26c0b18, 32'hc24eaed7} /* (8, 24, 15) {real, imag} */,
  {32'hc0eb1ba0, 32'hc16e0586} /* (8, 24, 14) {real, imag} */,
  {32'hc2b0074c, 32'hc2787344} /* (8, 24, 13) {real, imag} */,
  {32'hc2a91fba, 32'hc293f1ff} /* (8, 24, 12) {real, imag} */,
  {32'hc29c8a2b, 32'hc2236375} /* (8, 24, 11) {real, imag} */,
  {32'h40e21b00, 32'hc21ac8b2} /* (8, 24, 10) {real, imag} */,
  {32'h41df0b14, 32'h42c3e2ff} /* (8, 24, 9) {real, imag} */,
  {32'hc212654b, 32'hc2cdb43e} /* (8, 24, 8) {real, imag} */,
  {32'hc1d5d98a, 32'h428445f8} /* (8, 24, 7) {real, imag} */,
  {32'h4320199c, 32'hc1e4be22} /* (8, 24, 6) {real, imag} */,
  {32'hc362aa3a, 32'hc2df470a} /* (8, 24, 5) {real, imag} */,
  {32'h43101ed8, 32'hc2861a28} /* (8, 24, 4) {real, imag} */,
  {32'hc2c3779d, 32'h4291a886} /* (8, 24, 3) {real, imag} */,
  {32'hc4b7431a, 32'hc322aa0a} /* (8, 24, 2) {real, imag} */,
  {32'h456d9426, 32'h43c3ce30} /* (8, 24, 1) {real, imag} */,
  {32'h457d9060, 32'h00000000} /* (8, 24, 0) {real, imag} */,
  {32'h453f86a7, 32'hc39a5e50} /* (8, 23, 31) {real, imag} */,
  {32'hc4965d1b, 32'h43536c6a} /* (8, 23, 30) {real, imag} */,
  {32'hc33d6b04, 32'hc34f408f} /* (8, 23, 29) {real, imag} */,
  {32'h4323f0a0, 32'hc2266b3e} /* (8, 23, 28) {real, imag} */,
  {32'hc3aeab77, 32'h42b3c34e} /* (8, 23, 27) {real, imag} */,
  {32'hc0d40878, 32'hbf87c2a8} /* (8, 23, 26) {real, imag} */,
  {32'hc2018419, 32'hc2728cf9} /* (8, 23, 25) {real, imag} */,
  {32'hc2ca7b9f, 32'h41d813ca} /* (8, 23, 24) {real, imag} */,
  {32'h415ac8ee, 32'hc21e6d9f} /* (8, 23, 23) {real, imag} */,
  {32'hc279f0c2, 32'hc1af3978} /* (8, 23, 22) {real, imag} */,
  {32'hc006d3c0, 32'h42423347} /* (8, 23, 21) {real, imag} */,
  {32'hc2a21edc, 32'h412efd8e} /* (8, 23, 20) {real, imag} */,
  {32'hc0a584e4, 32'hc22c3626} /* (8, 23, 19) {real, imag} */,
  {32'h42ec5c23, 32'h423725e1} /* (8, 23, 18) {real, imag} */,
  {32'h424b559e, 32'h42bcffb6} /* (8, 23, 17) {real, imag} */,
  {32'hc2493156, 32'h00000000} /* (8, 23, 16) {real, imag} */,
  {32'h424b559e, 32'hc2bcffb6} /* (8, 23, 15) {real, imag} */,
  {32'h42ec5c23, 32'hc23725e1} /* (8, 23, 14) {real, imag} */,
  {32'hc0a584e4, 32'h422c3626} /* (8, 23, 13) {real, imag} */,
  {32'hc2a21edc, 32'hc12efd8e} /* (8, 23, 12) {real, imag} */,
  {32'hc006d3c0, 32'hc2423347} /* (8, 23, 11) {real, imag} */,
  {32'hc279f0c2, 32'h41af3978} /* (8, 23, 10) {real, imag} */,
  {32'h415ac8ee, 32'h421e6d9f} /* (8, 23, 9) {real, imag} */,
  {32'hc2ca7b9f, 32'hc1d813ca} /* (8, 23, 8) {real, imag} */,
  {32'hc2018419, 32'h42728cf9} /* (8, 23, 7) {real, imag} */,
  {32'hc0d40878, 32'h3f87c2a8} /* (8, 23, 6) {real, imag} */,
  {32'hc3aeab77, 32'hc2b3c34e} /* (8, 23, 5) {real, imag} */,
  {32'h4323f0a0, 32'h42266b3e} /* (8, 23, 4) {real, imag} */,
  {32'hc33d6b04, 32'h434f408f} /* (8, 23, 3) {real, imag} */,
  {32'hc4965d1b, 32'hc3536c6a} /* (8, 23, 2) {real, imag} */,
  {32'h453f86a7, 32'h439a5e50} /* (8, 23, 1) {real, imag} */,
  {32'h455029f0, 32'h00000000} /* (8, 23, 0) {real, imag} */,
  {32'h44f2dfe7, 32'hc38a0bee} /* (8, 22, 31) {real, imag} */,
  {32'hc45dce94, 32'h430a52dc} /* (8, 22, 30) {real, imag} */,
  {32'hc2228a52, 32'hc26e7806} /* (8, 22, 29) {real, imag} */,
  {32'h42d44344, 32'hc286a816} /* (8, 22, 28) {real, imag} */,
  {32'hc388edec, 32'h425a2813} /* (8, 22, 27) {real, imag} */,
  {32'h40a59012, 32'hc1130f04} /* (8, 22, 26) {real, imag} */,
  {32'hc2a83cb9, 32'h42090a9d} /* (8, 22, 25) {real, imag} */,
  {32'hc2b6871a, 32'h42209efc} /* (8, 22, 24) {real, imag} */,
  {32'hc199e9dd, 32'hc19a9dfd} /* (8, 22, 23) {real, imag} */,
  {32'h42aa5720, 32'h42729757} /* (8, 22, 22) {real, imag} */,
  {32'h42432115, 32'h42c4e3d3} /* (8, 22, 21) {real, imag} */,
  {32'h4234050a, 32'hc312a789} /* (8, 22, 20) {real, imag} */,
  {32'h42a07604, 32'hc1b5853e} /* (8, 22, 19) {real, imag} */,
  {32'hc1967d2a, 32'h41eb2d66} /* (8, 22, 18) {real, imag} */,
  {32'hc2907f48, 32'h3df29600} /* (8, 22, 17) {real, imag} */,
  {32'hc2b94f5a, 32'h00000000} /* (8, 22, 16) {real, imag} */,
  {32'hc2907f48, 32'hbdf29600} /* (8, 22, 15) {real, imag} */,
  {32'hc1967d2a, 32'hc1eb2d66} /* (8, 22, 14) {real, imag} */,
  {32'h42a07604, 32'h41b5853e} /* (8, 22, 13) {real, imag} */,
  {32'h4234050a, 32'h4312a789} /* (8, 22, 12) {real, imag} */,
  {32'h42432115, 32'hc2c4e3d3} /* (8, 22, 11) {real, imag} */,
  {32'h42aa5720, 32'hc2729757} /* (8, 22, 10) {real, imag} */,
  {32'hc199e9dd, 32'h419a9dfd} /* (8, 22, 9) {real, imag} */,
  {32'hc2b6871a, 32'hc2209efc} /* (8, 22, 8) {real, imag} */,
  {32'hc2a83cb9, 32'hc2090a9d} /* (8, 22, 7) {real, imag} */,
  {32'h40a59012, 32'h41130f04} /* (8, 22, 6) {real, imag} */,
  {32'hc388edec, 32'hc25a2813} /* (8, 22, 5) {real, imag} */,
  {32'h42d44344, 32'h4286a816} /* (8, 22, 4) {real, imag} */,
  {32'hc2228a52, 32'h426e7806} /* (8, 22, 3) {real, imag} */,
  {32'hc45dce94, 32'hc30a52dc} /* (8, 22, 2) {real, imag} */,
  {32'h44f2dfe7, 32'h438a0bee} /* (8, 22, 1) {real, imag} */,
  {32'h451792bc, 32'h00000000} /* (8, 22, 0) {real, imag} */,
  {32'h4405f0de, 32'hc286b03c} /* (8, 21, 31) {real, imag} */,
  {32'hc381fd60, 32'hc2d929df} /* (8, 21, 30) {real, imag} */,
  {32'h419b3e60, 32'hbfe14ca0} /* (8, 21, 29) {real, imag} */,
  {32'hc1f1efc8, 32'hc1a25594} /* (8, 21, 28) {real, imag} */,
  {32'hc2fb794d, 32'h41e617c9} /* (8, 21, 27) {real, imag} */,
  {32'h4193478b, 32'hc1e65904} /* (8, 21, 26) {real, imag} */,
  {32'hc2b940aa, 32'hc1dfb664} /* (8, 21, 25) {real, imag} */,
  {32'hc14184c0, 32'h42251674} /* (8, 21, 24) {real, imag} */,
  {32'hc1b70b0c, 32'hc27f0e8e} /* (8, 21, 23) {real, imag} */,
  {32'hc0e7ba70, 32'hc225104b} /* (8, 21, 22) {real, imag} */,
  {32'h422343c4, 32'h42abde5a} /* (8, 21, 21) {real, imag} */,
  {32'hc2524248, 32'hc209f6d6} /* (8, 21, 20) {real, imag} */,
  {32'h4266f966, 32'h42ded1c0} /* (8, 21, 19) {real, imag} */,
  {32'hc267093e, 32'h41b69c24} /* (8, 21, 18) {real, imag} */,
  {32'hc268c700, 32'h3f8e9600} /* (8, 21, 17) {real, imag} */,
  {32'hc282930a, 32'h00000000} /* (8, 21, 16) {real, imag} */,
  {32'hc268c700, 32'hbf8e9600} /* (8, 21, 15) {real, imag} */,
  {32'hc267093e, 32'hc1b69c24} /* (8, 21, 14) {real, imag} */,
  {32'h4266f966, 32'hc2ded1c0} /* (8, 21, 13) {real, imag} */,
  {32'hc2524248, 32'h4209f6d6} /* (8, 21, 12) {real, imag} */,
  {32'h422343c4, 32'hc2abde5a} /* (8, 21, 11) {real, imag} */,
  {32'hc0e7ba70, 32'h4225104b} /* (8, 21, 10) {real, imag} */,
  {32'hc1b70b0c, 32'h427f0e8e} /* (8, 21, 9) {real, imag} */,
  {32'hc14184c0, 32'hc2251674} /* (8, 21, 8) {real, imag} */,
  {32'hc2b940aa, 32'h41dfb664} /* (8, 21, 7) {real, imag} */,
  {32'h4193478b, 32'h41e65904} /* (8, 21, 6) {real, imag} */,
  {32'hc2fb794d, 32'hc1e617c9} /* (8, 21, 5) {real, imag} */,
  {32'hc1f1efc8, 32'h41a25594} /* (8, 21, 4) {real, imag} */,
  {32'h419b3e60, 32'h3fe14ca0} /* (8, 21, 3) {real, imag} */,
  {32'hc381fd60, 32'h42d929df} /* (8, 21, 2) {real, imag} */,
  {32'h4405f0de, 32'h4286b03c} /* (8, 21, 1) {real, imag} */,
  {32'h447ab9b4, 32'h00000000} /* (8, 21, 0) {real, imag} */,
  {32'hc4a34c60, 32'h41affb80} /* (8, 20, 31) {real, imag} */,
  {32'h440eea07, 32'hc3945a7a} /* (8, 20, 30) {real, imag} */,
  {32'hbfddfd80, 32'h421b33d9} /* (8, 20, 29) {real, imag} */,
  {32'hc2b4af84, 32'h427136a0} /* (8, 20, 28) {real, imag} */,
  {32'h428d4bd2, 32'hc270b464} /* (8, 20, 27) {real, imag} */,
  {32'h4188e11f, 32'h427ad1e0} /* (8, 20, 26) {real, imag} */,
  {32'hc1e82178, 32'h403134b0} /* (8, 20, 25) {real, imag} */,
  {32'h427237fa, 32'h42094aac} /* (8, 20, 24) {real, imag} */,
  {32'h424ddb83, 32'hc2d3595f} /* (8, 20, 23) {real, imag} */,
  {32'h42ac1b22, 32'hc304b744} /* (8, 20, 22) {real, imag} */,
  {32'h428701fe, 32'hc28bdbdc} /* (8, 20, 21) {real, imag} */,
  {32'hbffd6650, 32'h40a64bc2} /* (8, 20, 20) {real, imag} */,
  {32'hc19b0e97, 32'h412317f4} /* (8, 20, 19) {real, imag} */,
  {32'hc260c151, 32'hc11fcf5c} /* (8, 20, 18) {real, imag} */,
  {32'h411428f8, 32'h41d21a66} /* (8, 20, 17) {real, imag} */,
  {32'hc29e21b3, 32'h00000000} /* (8, 20, 16) {real, imag} */,
  {32'h411428f8, 32'hc1d21a66} /* (8, 20, 15) {real, imag} */,
  {32'hc260c151, 32'h411fcf5c} /* (8, 20, 14) {real, imag} */,
  {32'hc19b0e97, 32'hc12317f4} /* (8, 20, 13) {real, imag} */,
  {32'hbffd6650, 32'hc0a64bc2} /* (8, 20, 12) {real, imag} */,
  {32'h428701fe, 32'h428bdbdc} /* (8, 20, 11) {real, imag} */,
  {32'h42ac1b22, 32'h4304b744} /* (8, 20, 10) {real, imag} */,
  {32'h424ddb83, 32'h42d3595f} /* (8, 20, 9) {real, imag} */,
  {32'h427237fa, 32'hc2094aac} /* (8, 20, 8) {real, imag} */,
  {32'hc1e82178, 32'hc03134b0} /* (8, 20, 7) {real, imag} */,
  {32'h4188e11f, 32'hc27ad1e0} /* (8, 20, 6) {real, imag} */,
  {32'h428d4bd2, 32'h4270b464} /* (8, 20, 5) {real, imag} */,
  {32'hc2b4af84, 32'hc27136a0} /* (8, 20, 4) {real, imag} */,
  {32'hbfddfd80, 32'hc21b33d9} /* (8, 20, 3) {real, imag} */,
  {32'h440eea07, 32'h43945a7a} /* (8, 20, 2) {real, imag} */,
  {32'hc4a34c60, 32'hc1affb80} /* (8, 20, 1) {real, imag} */,
  {32'hc4018449, 32'h00000000} /* (8, 20, 0) {real, imag} */,
  {32'hc51ed520, 32'h4208f0d0} /* (8, 19, 31) {real, imag} */,
  {32'h4485f5cf, 32'hc38bc138} /* (8, 19, 30) {real, imag} */,
  {32'h412af2c4, 32'h41f9035c} /* (8, 19, 29) {real, imag} */,
  {32'hc365cfd4, 32'hc3040507} /* (8, 19, 28) {real, imag} */,
  {32'h438209fd, 32'hc2f4d9f5} /* (8, 19, 27) {real, imag} */,
  {32'h42bd0016, 32'hc1f7bacf} /* (8, 19, 26) {real, imag} */,
  {32'h42457aa4, 32'h430fca82} /* (8, 19, 25) {real, imag} */,
  {32'h41350af8, 32'hc21acf42} /* (8, 19, 24) {real, imag} */,
  {32'hc281a2e2, 32'hc295e9f8} /* (8, 19, 23) {real, imag} */,
  {32'h42063657, 32'h43336a9b} /* (8, 19, 22) {real, imag} */,
  {32'hc2f8d02c, 32'hc1b9aa5c} /* (8, 19, 21) {real, imag} */,
  {32'h41f0407c, 32'hc139bbab} /* (8, 19, 20) {real, imag} */,
  {32'h42ca2482, 32'h42294082} /* (8, 19, 19) {real, imag} */,
  {32'hc2c67553, 32'hc273e9d0} /* (8, 19, 18) {real, imag} */,
  {32'h41e5bfb0, 32'hc15bb05a} /* (8, 19, 17) {real, imag} */,
  {32'hc0f9d920, 32'h00000000} /* (8, 19, 16) {real, imag} */,
  {32'h41e5bfb0, 32'h415bb05a} /* (8, 19, 15) {real, imag} */,
  {32'hc2c67553, 32'h4273e9d0} /* (8, 19, 14) {real, imag} */,
  {32'h42ca2482, 32'hc2294082} /* (8, 19, 13) {real, imag} */,
  {32'h41f0407c, 32'h4139bbab} /* (8, 19, 12) {real, imag} */,
  {32'hc2f8d02c, 32'h41b9aa5c} /* (8, 19, 11) {real, imag} */,
  {32'h42063657, 32'hc3336a9b} /* (8, 19, 10) {real, imag} */,
  {32'hc281a2e2, 32'h4295e9f8} /* (8, 19, 9) {real, imag} */,
  {32'h41350af8, 32'h421acf42} /* (8, 19, 8) {real, imag} */,
  {32'h42457aa4, 32'hc30fca82} /* (8, 19, 7) {real, imag} */,
  {32'h42bd0016, 32'h41f7bacf} /* (8, 19, 6) {real, imag} */,
  {32'h438209fd, 32'h42f4d9f5} /* (8, 19, 5) {real, imag} */,
  {32'hc365cfd4, 32'h43040507} /* (8, 19, 4) {real, imag} */,
  {32'h412af2c4, 32'hc1f9035c} /* (8, 19, 3) {real, imag} */,
  {32'h4485f5cf, 32'h438bc138} /* (8, 19, 2) {real, imag} */,
  {32'hc51ed520, 32'hc208f0d0} /* (8, 19, 1) {real, imag} */,
  {32'hc4b7bdc0, 32'h00000000} /* (8, 19, 0) {real, imag} */,
  {32'hc5579699, 32'h43878570} /* (8, 18, 31) {real, imag} */,
  {32'h449ee1d2, 32'hc38db865} /* (8, 18, 30) {real, imag} */,
  {32'hc3190cfe, 32'hc2e475e3} /* (8, 18, 29) {real, imag} */,
  {32'hc3a72d34, 32'hc26841af} /* (8, 18, 28) {real, imag} */,
  {32'h43832f86, 32'h428e0b5c} /* (8, 18, 27) {real, imag} */,
  {32'h426b41f6, 32'hc2c7c270} /* (8, 18, 26) {real, imag} */,
  {32'hc05978c8, 32'h42ba53d6} /* (8, 18, 25) {real, imag} */,
  {32'h431f32f2, 32'h42814065} /* (8, 18, 24) {real, imag} */,
  {32'hc200a6d4, 32'h421d6c46} /* (8, 18, 23) {real, imag} */,
  {32'hc213eae4, 32'hc29c30a3} /* (8, 18, 22) {real, imag} */,
  {32'h423e2998, 32'hc244b0a1} /* (8, 18, 21) {real, imag} */,
  {32'hc237540e, 32'h4208d3e8} /* (8, 18, 20) {real, imag} */,
  {32'hc0dc9f34, 32'hc2c8f57a} /* (8, 18, 19) {real, imag} */,
  {32'h4260a8a0, 32'hc1e9acf6} /* (8, 18, 18) {real, imag} */,
  {32'hc10e23a4, 32'h41cbf776} /* (8, 18, 17) {real, imag} */,
  {32'h4088b3ae, 32'h00000000} /* (8, 18, 16) {real, imag} */,
  {32'hc10e23a4, 32'hc1cbf776} /* (8, 18, 15) {real, imag} */,
  {32'h4260a8a0, 32'h41e9acf6} /* (8, 18, 14) {real, imag} */,
  {32'hc0dc9f34, 32'h42c8f57a} /* (8, 18, 13) {real, imag} */,
  {32'hc237540e, 32'hc208d3e8} /* (8, 18, 12) {real, imag} */,
  {32'h423e2998, 32'h4244b0a1} /* (8, 18, 11) {real, imag} */,
  {32'hc213eae4, 32'h429c30a3} /* (8, 18, 10) {real, imag} */,
  {32'hc200a6d4, 32'hc21d6c46} /* (8, 18, 9) {real, imag} */,
  {32'h431f32f2, 32'hc2814065} /* (8, 18, 8) {real, imag} */,
  {32'hc05978c8, 32'hc2ba53d6} /* (8, 18, 7) {real, imag} */,
  {32'h426b41f6, 32'h42c7c270} /* (8, 18, 6) {real, imag} */,
  {32'h43832f86, 32'hc28e0b5c} /* (8, 18, 5) {real, imag} */,
  {32'hc3a72d34, 32'h426841af} /* (8, 18, 4) {real, imag} */,
  {32'hc3190cfe, 32'h42e475e3} /* (8, 18, 3) {real, imag} */,
  {32'h449ee1d2, 32'h438db865} /* (8, 18, 2) {real, imag} */,
  {32'hc5579699, 32'hc3878570} /* (8, 18, 1) {real, imag} */,
  {32'hc50e7556, 32'h00000000} /* (8, 18, 0) {real, imag} */,
  {32'hc571653b, 32'h438f8c82} /* (8, 17, 31) {real, imag} */,
  {32'h449fcc1b, 32'hc34fb7cc} /* (8, 17, 30) {real, imag} */,
  {32'hc240b305, 32'hc24e54db} /* (8, 17, 29) {real, imag} */,
  {32'hc3003335, 32'h42ac0ae9} /* (8, 17, 28) {real, imag} */,
  {32'h4389ea8e, 32'h43013104} /* (8, 17, 27) {real, imag} */,
  {32'h43654d4a, 32'hc297b235} /* (8, 17, 26) {real, imag} */,
  {32'hc2066266, 32'h413476e6} /* (8, 17, 25) {real, imag} */,
  {32'h42a29442, 32'h42eea609} /* (8, 17, 24) {real, imag} */,
  {32'h429b117f, 32'hc22d5714} /* (8, 17, 23) {real, imag} */,
  {32'h41883e7c, 32'hc24c013d} /* (8, 17, 22) {real, imag} */,
  {32'hc20cabcd, 32'hc1bfc788} /* (8, 17, 21) {real, imag} */,
  {32'hc0cd283e, 32'hc2a3dc1b} /* (8, 17, 20) {real, imag} */,
  {32'hc1b87d95, 32'hc2b7cfd8} /* (8, 17, 19) {real, imag} */,
  {32'h4244dbc2, 32'hc1c6d26e} /* (8, 17, 18) {real, imag} */,
  {32'hc20210be, 32'h42183892} /* (8, 17, 17) {real, imag} */,
  {32'h41b0330e, 32'h00000000} /* (8, 17, 16) {real, imag} */,
  {32'hc20210be, 32'hc2183892} /* (8, 17, 15) {real, imag} */,
  {32'h4244dbc2, 32'h41c6d26e} /* (8, 17, 14) {real, imag} */,
  {32'hc1b87d95, 32'h42b7cfd8} /* (8, 17, 13) {real, imag} */,
  {32'hc0cd283e, 32'h42a3dc1b} /* (8, 17, 12) {real, imag} */,
  {32'hc20cabcd, 32'h41bfc788} /* (8, 17, 11) {real, imag} */,
  {32'h41883e7c, 32'h424c013d} /* (8, 17, 10) {real, imag} */,
  {32'h429b117f, 32'h422d5714} /* (8, 17, 9) {real, imag} */,
  {32'h42a29442, 32'hc2eea609} /* (8, 17, 8) {real, imag} */,
  {32'hc2066266, 32'hc13476e6} /* (8, 17, 7) {real, imag} */,
  {32'h43654d4a, 32'h4297b235} /* (8, 17, 6) {real, imag} */,
  {32'h4389ea8e, 32'hc3013104} /* (8, 17, 5) {real, imag} */,
  {32'hc3003335, 32'hc2ac0ae9} /* (8, 17, 4) {real, imag} */,
  {32'hc240b305, 32'h424e54db} /* (8, 17, 3) {real, imag} */,
  {32'h449fcc1b, 32'h434fb7cc} /* (8, 17, 2) {real, imag} */,
  {32'hc571653b, 32'hc38f8c82} /* (8, 17, 1) {real, imag} */,
  {32'hc5425110, 32'h00000000} /* (8, 17, 0) {real, imag} */,
  {32'hc5811c96, 32'h43886fac} /* (8, 16, 31) {real, imag} */,
  {32'h44a9c94a, 32'hc378ac38} /* (8, 16, 30) {real, imag} */,
  {32'hc29d1317, 32'hc1f5597a} /* (8, 16, 29) {real, imag} */,
  {32'hc2f68f38, 32'h416c4778} /* (8, 16, 28) {real, imag} */,
  {32'h438d6641, 32'hc1d2e4c4} /* (8, 16, 27) {real, imag} */,
  {32'h42b40e88, 32'hc1da9e40} /* (8, 16, 26) {real, imag} */,
  {32'hc03ed030, 32'h42037256} /* (8, 16, 25) {real, imag} */,
  {32'h42460e9c, 32'h40fa766a} /* (8, 16, 24) {real, imag} */,
  {32'h42b72d22, 32'hc1ced608} /* (8, 16, 23) {real, imag} */,
  {32'h42749520, 32'hc109e570} /* (8, 16, 22) {real, imag} */,
  {32'h425ca64b, 32'hc1fd2f61} /* (8, 16, 21) {real, imag} */,
  {32'hc1ab1208, 32'hc3030d39} /* (8, 16, 20) {real, imag} */,
  {32'h425bbb82, 32'hc2021b83} /* (8, 16, 19) {real, imag} */,
  {32'hc260f8d9, 32'hc1a4bc00} /* (8, 16, 18) {real, imag} */,
  {32'h417c8118, 32'h421372fa} /* (8, 16, 17) {real, imag} */,
  {32'hc246b56b, 32'h00000000} /* (8, 16, 16) {real, imag} */,
  {32'h417c8118, 32'hc21372fa} /* (8, 16, 15) {real, imag} */,
  {32'hc260f8d9, 32'h41a4bc00} /* (8, 16, 14) {real, imag} */,
  {32'h425bbb82, 32'h42021b83} /* (8, 16, 13) {real, imag} */,
  {32'hc1ab1208, 32'h43030d39} /* (8, 16, 12) {real, imag} */,
  {32'h425ca64b, 32'h41fd2f61} /* (8, 16, 11) {real, imag} */,
  {32'h42749520, 32'h4109e570} /* (8, 16, 10) {real, imag} */,
  {32'h42b72d22, 32'h41ced608} /* (8, 16, 9) {real, imag} */,
  {32'h42460e9c, 32'hc0fa766a} /* (8, 16, 8) {real, imag} */,
  {32'hc03ed030, 32'hc2037256} /* (8, 16, 7) {real, imag} */,
  {32'h42b40e88, 32'h41da9e40} /* (8, 16, 6) {real, imag} */,
  {32'h438d6641, 32'h41d2e4c4} /* (8, 16, 5) {real, imag} */,
  {32'hc2f68f38, 32'hc16c4778} /* (8, 16, 4) {real, imag} */,
  {32'hc29d1317, 32'h41f5597a} /* (8, 16, 3) {real, imag} */,
  {32'h44a9c94a, 32'h4378ac38} /* (8, 16, 2) {real, imag} */,
  {32'hc5811c96, 32'hc3886fac} /* (8, 16, 1) {real, imag} */,
  {32'hc5409f22, 32'h00000000} /* (8, 16, 0) {real, imag} */,
  {32'hc580454e, 32'h437d90bc} /* (8, 15, 31) {real, imag} */,
  {32'h44b2f205, 32'hc350d6f0} /* (8, 15, 30) {real, imag} */,
  {32'hc1cfc082, 32'h4295221a} /* (8, 15, 29) {real, imag} */,
  {32'hc372be83, 32'h42ac21cf} /* (8, 15, 28) {real, imag} */,
  {32'h431f3267, 32'hc0fa0a70} /* (8, 15, 27) {real, imag} */,
  {32'h433097d2, 32'h3f23dd80} /* (8, 15, 26) {real, imag} */,
  {32'h42bb905f, 32'hc27d819c} /* (8, 15, 25) {real, imag} */,
  {32'h42b0e452, 32'h42abdd71} /* (8, 15, 24) {real, imag} */,
  {32'hc15ba306, 32'hc1836ae3} /* (8, 15, 23) {real, imag} */,
  {32'hc248b4fa, 32'hc1925292} /* (8, 15, 22) {real, imag} */,
  {32'h427ecdf1, 32'hc28e622e} /* (8, 15, 21) {real, imag} */,
  {32'hc1880e70, 32'h42646a86} /* (8, 15, 20) {real, imag} */,
  {32'h41a30c23, 32'h428f98f4} /* (8, 15, 19) {real, imag} */,
  {32'h422adcc6, 32'hc2425131} /* (8, 15, 18) {real, imag} */,
  {32'hc1e3287b, 32'hc0571618} /* (8, 15, 17) {real, imag} */,
  {32'hbf2f8f00, 32'h00000000} /* (8, 15, 16) {real, imag} */,
  {32'hc1e3287b, 32'h40571618} /* (8, 15, 15) {real, imag} */,
  {32'h422adcc6, 32'h42425131} /* (8, 15, 14) {real, imag} */,
  {32'h41a30c23, 32'hc28f98f4} /* (8, 15, 13) {real, imag} */,
  {32'hc1880e70, 32'hc2646a86} /* (8, 15, 12) {real, imag} */,
  {32'h427ecdf1, 32'h428e622e} /* (8, 15, 11) {real, imag} */,
  {32'hc248b4fa, 32'h41925292} /* (8, 15, 10) {real, imag} */,
  {32'hc15ba306, 32'h41836ae3} /* (8, 15, 9) {real, imag} */,
  {32'h42b0e452, 32'hc2abdd71} /* (8, 15, 8) {real, imag} */,
  {32'h42bb905f, 32'h427d819c} /* (8, 15, 7) {real, imag} */,
  {32'h433097d2, 32'hbf23dd80} /* (8, 15, 6) {real, imag} */,
  {32'h431f3267, 32'h40fa0a70} /* (8, 15, 5) {real, imag} */,
  {32'hc372be83, 32'hc2ac21cf} /* (8, 15, 4) {real, imag} */,
  {32'hc1cfc082, 32'hc295221a} /* (8, 15, 3) {real, imag} */,
  {32'h44b2f205, 32'h4350d6f0} /* (8, 15, 2) {real, imag} */,
  {32'hc580454e, 32'hc37d90bc} /* (8, 15, 1) {real, imag} */,
  {32'hc53a4a9c, 32'h00000000} /* (8, 15, 0) {real, imag} */,
  {32'hc55d6df3, 32'h4368b670} /* (8, 14, 31) {real, imag} */,
  {32'h44ac3086, 32'hc36beda2} /* (8, 14, 30) {real, imag} */,
  {32'h4264d451, 32'h421de046} /* (8, 14, 29) {real, imag} */,
  {32'hc38c91e0, 32'h4223a5d3} /* (8, 14, 28) {real, imag} */,
  {32'h42a9658a, 32'hc371507c} /* (8, 14, 27) {real, imag} */,
  {32'h4247a3f2, 32'hc229a2b0} /* (8, 14, 26) {real, imag} */,
  {32'hc0d12b04, 32'h4291fe7e} /* (8, 14, 25) {real, imag} */,
  {32'h41426fa0, 32'hc196a348} /* (8, 14, 24) {real, imag} */,
  {32'hc1f6b77b, 32'hc2dff245} /* (8, 14, 23) {real, imag} */,
  {32'hc28722e4, 32'h42824e55} /* (8, 14, 22) {real, imag} */,
  {32'h42196234, 32'hc212aaa3} /* (8, 14, 21) {real, imag} */,
  {32'h4241930a, 32'hc2894843} /* (8, 14, 20) {real, imag} */,
  {32'hc1816407, 32'hc0db3de0} /* (8, 14, 19) {real, imag} */,
  {32'hc28db9e7, 32'hc1f4b7ba} /* (8, 14, 18) {real, imag} */,
  {32'hc12621b0, 32'hc0b30ad8} /* (8, 14, 17) {real, imag} */,
  {32'hc1a0b2c2, 32'h00000000} /* (8, 14, 16) {real, imag} */,
  {32'hc12621b0, 32'h40b30ad8} /* (8, 14, 15) {real, imag} */,
  {32'hc28db9e7, 32'h41f4b7ba} /* (8, 14, 14) {real, imag} */,
  {32'hc1816407, 32'h40db3de0} /* (8, 14, 13) {real, imag} */,
  {32'h4241930a, 32'h42894843} /* (8, 14, 12) {real, imag} */,
  {32'h42196234, 32'h4212aaa3} /* (8, 14, 11) {real, imag} */,
  {32'hc28722e4, 32'hc2824e55} /* (8, 14, 10) {real, imag} */,
  {32'hc1f6b77b, 32'h42dff245} /* (8, 14, 9) {real, imag} */,
  {32'h41426fa0, 32'h4196a348} /* (8, 14, 8) {real, imag} */,
  {32'hc0d12b04, 32'hc291fe7e} /* (8, 14, 7) {real, imag} */,
  {32'h4247a3f2, 32'h4229a2b0} /* (8, 14, 6) {real, imag} */,
  {32'h42a9658a, 32'h4371507c} /* (8, 14, 5) {real, imag} */,
  {32'hc38c91e0, 32'hc223a5d3} /* (8, 14, 4) {real, imag} */,
  {32'h4264d451, 32'hc21de046} /* (8, 14, 3) {real, imag} */,
  {32'h44ac3086, 32'h436beda2} /* (8, 14, 2) {real, imag} */,
  {32'hc55d6df3, 32'hc368b670} /* (8, 14, 1) {real, imag} */,
  {32'hc539979a, 32'h00000000} /* (8, 14, 0) {real, imag} */,
  {32'hc53ebcd2, 32'h42ebc4f8} /* (8, 13, 31) {real, imag} */,
  {32'h449b1285, 32'hc39d436e} /* (8, 13, 30) {real, imag} */,
  {32'h428ce678, 32'h421fa31a} /* (8, 13, 29) {real, imag} */,
  {32'hc350a666, 32'h4254890c} /* (8, 13, 28) {real, imag} */,
  {32'h42f44dad, 32'hc2f545cd} /* (8, 13, 27) {real, imag} */,
  {32'hc208f5e8, 32'hc1975e9f} /* (8, 13, 26) {real, imag} */,
  {32'hc31fea79, 32'h42055f43} /* (8, 13, 25) {real, imag} */,
  {32'h4342b19e, 32'hc308451c} /* (8, 13, 24) {real, imag} */,
  {32'h4252ec00, 32'hc1357d0c} /* (8, 13, 23) {real, imag} */,
  {32'h425db003, 32'h4205d38c} /* (8, 13, 22) {real, imag} */,
  {32'h42ac2ad8, 32'hc22269d4} /* (8, 13, 21) {real, imag} */,
  {32'hc274b2bc, 32'hc1cfeb82} /* (8, 13, 20) {real, imag} */,
  {32'hc14f22a0, 32'h41af514c} /* (8, 13, 19) {real, imag} */,
  {32'h42157ed2, 32'hc203d4fe} /* (8, 13, 18) {real, imag} */,
  {32'h400d499c, 32'h3f8368d0} /* (8, 13, 17) {real, imag} */,
  {32'hc2638cf8, 32'h00000000} /* (8, 13, 16) {real, imag} */,
  {32'h400d499c, 32'hbf8368d0} /* (8, 13, 15) {real, imag} */,
  {32'h42157ed2, 32'h4203d4fe} /* (8, 13, 14) {real, imag} */,
  {32'hc14f22a0, 32'hc1af514c} /* (8, 13, 13) {real, imag} */,
  {32'hc274b2bc, 32'h41cfeb82} /* (8, 13, 12) {real, imag} */,
  {32'h42ac2ad8, 32'h422269d4} /* (8, 13, 11) {real, imag} */,
  {32'h425db003, 32'hc205d38c} /* (8, 13, 10) {real, imag} */,
  {32'h4252ec00, 32'h41357d0c} /* (8, 13, 9) {real, imag} */,
  {32'h4342b19e, 32'h4308451c} /* (8, 13, 8) {real, imag} */,
  {32'hc31fea79, 32'hc2055f43} /* (8, 13, 7) {real, imag} */,
  {32'hc208f5e8, 32'h41975e9f} /* (8, 13, 6) {real, imag} */,
  {32'h42f44dad, 32'h42f545cd} /* (8, 13, 5) {real, imag} */,
  {32'hc350a666, 32'hc254890c} /* (8, 13, 4) {real, imag} */,
  {32'h428ce678, 32'hc21fa31a} /* (8, 13, 3) {real, imag} */,
  {32'h449b1285, 32'h439d436e} /* (8, 13, 2) {real, imag} */,
  {32'hc53ebcd2, 32'hc2ebc4f8} /* (8, 13, 1) {real, imag} */,
  {32'hc5126c5e, 32'h00000000} /* (8, 13, 0) {real, imag} */,
  {32'hc50a6992, 32'hc2a0b9c0} /* (8, 12, 31) {real, imag} */,
  {32'h44835d8c, 32'hc1dddec8} /* (8, 12, 30) {real, imag} */,
  {32'h435e046c, 32'h4109a210} /* (8, 12, 29) {real, imag} */,
  {32'hc2825480, 32'hc30cb669} /* (8, 12, 28) {real, imag} */,
  {32'h42f1625a, 32'hc24e6cac} /* (8, 12, 27) {real, imag} */,
  {32'h42946556, 32'hc21095e8} /* (8, 12, 26) {real, imag} */,
  {32'hc307d481, 32'h4256f749} /* (8, 12, 25) {real, imag} */,
  {32'h4222d340, 32'hc288b8e3} /* (8, 12, 24) {real, imag} */,
  {32'hc20d145f, 32'h4254e256} /* (8, 12, 23) {real, imag} */,
  {32'hc2642af4, 32'h42c362c4} /* (8, 12, 22) {real, imag} */,
  {32'hc04e3a90, 32'hc2581d1e} /* (8, 12, 21) {real, imag} */,
  {32'hc1a86ff3, 32'hc1ffdbc4} /* (8, 12, 20) {real, imag} */,
  {32'h4280116c, 32'h4087b114} /* (8, 12, 19) {real, imag} */,
  {32'hc28ae7de, 32'hc26e8f3b} /* (8, 12, 18) {real, imag} */,
  {32'hbfc0ec40, 32'hc1174f10} /* (8, 12, 17) {real, imag} */,
  {32'h403f5a80, 32'h00000000} /* (8, 12, 16) {real, imag} */,
  {32'hbfc0ec40, 32'h41174f10} /* (8, 12, 15) {real, imag} */,
  {32'hc28ae7de, 32'h426e8f3b} /* (8, 12, 14) {real, imag} */,
  {32'h4280116c, 32'hc087b114} /* (8, 12, 13) {real, imag} */,
  {32'hc1a86ff3, 32'h41ffdbc4} /* (8, 12, 12) {real, imag} */,
  {32'hc04e3a90, 32'h42581d1e} /* (8, 12, 11) {real, imag} */,
  {32'hc2642af4, 32'hc2c362c4} /* (8, 12, 10) {real, imag} */,
  {32'hc20d145f, 32'hc254e256} /* (8, 12, 9) {real, imag} */,
  {32'h4222d340, 32'h4288b8e3} /* (8, 12, 8) {real, imag} */,
  {32'hc307d481, 32'hc256f749} /* (8, 12, 7) {real, imag} */,
  {32'h42946556, 32'h421095e8} /* (8, 12, 6) {real, imag} */,
  {32'h42f1625a, 32'h424e6cac} /* (8, 12, 5) {real, imag} */,
  {32'hc2825480, 32'h430cb669} /* (8, 12, 4) {real, imag} */,
  {32'h435e046c, 32'hc109a210} /* (8, 12, 3) {real, imag} */,
  {32'h44835d8c, 32'h41dddec8} /* (8, 12, 2) {real, imag} */,
  {32'hc50a6992, 32'h42a0b9c0} /* (8, 12, 1) {real, imag} */,
  {32'hc4c2b7bc, 32'h00000000} /* (8, 12, 0) {real, imag} */,
  {32'hc48464ef, 32'hc392aaf1} /* (8, 11, 31) {real, imag} */,
  {32'h4405441e, 32'h416e43b8} /* (8, 11, 30) {real, imag} */,
  {32'h4350db9c, 32'h42995d98} /* (8, 11, 29) {real, imag} */,
  {32'hc318f5bd, 32'hc3329e7a} /* (8, 11, 28) {real, imag} */,
  {32'h40f190f0, 32'hc29e444a} /* (8, 11, 27) {real, imag} */,
  {32'h41da9917, 32'hc2d6f2c7} /* (8, 11, 26) {real, imag} */,
  {32'hc30980cd, 32'hc321e178} /* (8, 11, 25) {real, imag} */,
  {32'hc11099f0, 32'hc2f24d0e} /* (8, 11, 24) {real, imag} */,
  {32'h42b010e9, 32'h42640bbe} /* (8, 11, 23) {real, imag} */,
  {32'h42cc92ef, 32'h4250b86b} /* (8, 11, 22) {real, imag} */,
  {32'hc19ea28f, 32'hc14f1948} /* (8, 11, 21) {real, imag} */,
  {32'h40519000, 32'hc22d2436} /* (8, 11, 20) {real, imag} */,
  {32'hc260e786, 32'h41ab9788} /* (8, 11, 19) {real, imag} */,
  {32'h422ef5d2, 32'hc2426368} /* (8, 11, 18) {real, imag} */,
  {32'h41da2d9b, 32'hc08428f0} /* (8, 11, 17) {real, imag} */,
  {32'hc2a7ea3c, 32'h00000000} /* (8, 11, 16) {real, imag} */,
  {32'h41da2d9b, 32'h408428f0} /* (8, 11, 15) {real, imag} */,
  {32'h422ef5d2, 32'h42426368} /* (8, 11, 14) {real, imag} */,
  {32'hc260e786, 32'hc1ab9788} /* (8, 11, 13) {real, imag} */,
  {32'h40519000, 32'h422d2436} /* (8, 11, 12) {real, imag} */,
  {32'hc19ea28f, 32'h414f1948} /* (8, 11, 11) {real, imag} */,
  {32'h42cc92ef, 32'hc250b86b} /* (8, 11, 10) {real, imag} */,
  {32'h42b010e9, 32'hc2640bbe} /* (8, 11, 9) {real, imag} */,
  {32'hc11099f0, 32'h42f24d0e} /* (8, 11, 8) {real, imag} */,
  {32'hc30980cd, 32'h4321e178} /* (8, 11, 7) {real, imag} */,
  {32'h41da9917, 32'h42d6f2c7} /* (8, 11, 6) {real, imag} */,
  {32'h40f190f0, 32'h429e444a} /* (8, 11, 5) {real, imag} */,
  {32'hc318f5bd, 32'h43329e7a} /* (8, 11, 4) {real, imag} */,
  {32'h4350db9c, 32'hc2995d98} /* (8, 11, 3) {real, imag} */,
  {32'h4405441e, 32'hc16e43b8} /* (8, 11, 2) {real, imag} */,
  {32'hc48464ef, 32'h4392aaf1} /* (8, 11, 1) {real, imag} */,
  {32'hc41bb374, 32'h00000000} /* (8, 11, 0) {real, imag} */,
  {32'h440b928a, 32'hc42ea12a} /* (8, 10, 31) {real, imag} */,
  {32'hc38df841, 32'h4346f7c4} /* (8, 10, 30) {real, imag} */,
  {32'h42e3e56b, 32'h423a578a} /* (8, 10, 29) {real, imag} */,
  {32'hc25e8920, 32'hc32be61f} /* (8, 10, 28) {real, imag} */,
  {32'hc2e9966a, 32'h43179a77} /* (8, 10, 27) {real, imag} */,
  {32'hc0b42f72, 32'hc1a3c336} /* (8, 10, 26) {real, imag} */,
  {32'h41b53f08, 32'hc30a3e6b} /* (8, 10, 25) {real, imag} */,
  {32'h42b2c1b6, 32'hc2d1224a} /* (8, 10, 24) {real, imag} */,
  {32'hc20b3a12, 32'hc186e6b9} /* (8, 10, 23) {real, imag} */,
  {32'h42765901, 32'h428e588e} /* (8, 10, 22) {real, imag} */,
  {32'h4021b4c0, 32'h41f4542c} /* (8, 10, 21) {real, imag} */,
  {32'hc254ce52, 32'h4230abdc} /* (8, 10, 20) {real, imag} */,
  {32'hbfb116a0, 32'h42b5a9a2} /* (8, 10, 19) {real, imag} */,
  {32'h428a8e8a, 32'h41e01086} /* (8, 10, 18) {real, imag} */,
  {32'hc11192ee, 32'hc29faf14} /* (8, 10, 17) {real, imag} */,
  {32'hc0c0a2f8, 32'h00000000} /* (8, 10, 16) {real, imag} */,
  {32'hc11192ee, 32'h429faf14} /* (8, 10, 15) {real, imag} */,
  {32'h428a8e8a, 32'hc1e01086} /* (8, 10, 14) {real, imag} */,
  {32'hbfb116a0, 32'hc2b5a9a2} /* (8, 10, 13) {real, imag} */,
  {32'hc254ce52, 32'hc230abdc} /* (8, 10, 12) {real, imag} */,
  {32'h4021b4c0, 32'hc1f4542c} /* (8, 10, 11) {real, imag} */,
  {32'h42765901, 32'hc28e588e} /* (8, 10, 10) {real, imag} */,
  {32'hc20b3a12, 32'h4186e6b9} /* (8, 10, 9) {real, imag} */,
  {32'h42b2c1b6, 32'h42d1224a} /* (8, 10, 8) {real, imag} */,
  {32'h41b53f08, 32'h430a3e6b} /* (8, 10, 7) {real, imag} */,
  {32'hc0b42f72, 32'h41a3c336} /* (8, 10, 6) {real, imag} */,
  {32'hc2e9966a, 32'hc3179a77} /* (8, 10, 5) {real, imag} */,
  {32'hc25e8920, 32'h432be61f} /* (8, 10, 4) {real, imag} */,
  {32'h42e3e56b, 32'hc23a578a} /* (8, 10, 3) {real, imag} */,
  {32'hc38df841, 32'hc346f7c4} /* (8, 10, 2) {real, imag} */,
  {32'h440b928a, 32'h442ea12a} /* (8, 10, 1) {real, imag} */,
  {32'h4472eb51, 32'h00000000} /* (8, 10, 0) {real, imag} */,
  {32'h44f30a1e, 32'hc47e1134} /* (8, 9, 31) {real, imag} */,
  {32'hc448360a, 32'h43e03f2d} /* (8, 9, 30) {real, imag} */,
  {32'h4240d132, 32'hc3125491} /* (8, 9, 29) {real, imag} */,
  {32'h43087d6a, 32'hc2d388db} /* (8, 9, 28) {real, imag} */,
  {32'hc32cc492, 32'h42ae83ea} /* (8, 9, 27) {real, imag} */,
  {32'h427db2c1, 32'h41098261} /* (8, 9, 26) {real, imag} */,
  {32'hc26e9df5, 32'h4233ad71} /* (8, 9, 25) {real, imag} */,
  {32'h42c595b1, 32'h41bb661e} /* (8, 9, 24) {real, imag} */,
  {32'h42845f5d, 32'h4231de7f} /* (8, 9, 23) {real, imag} */,
  {32'hc297d28b, 32'h425409e0} /* (8, 9, 22) {real, imag} */,
  {32'h42492d84, 32'hc2b97c72} /* (8, 9, 21) {real, imag} */,
  {32'hc21dfd75, 32'h4271ded4} /* (8, 9, 20) {real, imag} */,
  {32'h42544936, 32'hc25a9da6} /* (8, 9, 19) {real, imag} */,
  {32'h429e2af1, 32'h4075f770} /* (8, 9, 18) {real, imag} */,
  {32'hc246f674, 32'hc1067604} /* (8, 9, 17) {real, imag} */,
  {32'hc1a5cfc0, 32'h00000000} /* (8, 9, 16) {real, imag} */,
  {32'hc246f674, 32'h41067604} /* (8, 9, 15) {real, imag} */,
  {32'h429e2af1, 32'hc075f770} /* (8, 9, 14) {real, imag} */,
  {32'h42544936, 32'h425a9da6} /* (8, 9, 13) {real, imag} */,
  {32'hc21dfd75, 32'hc271ded4} /* (8, 9, 12) {real, imag} */,
  {32'h42492d84, 32'h42b97c72} /* (8, 9, 11) {real, imag} */,
  {32'hc297d28b, 32'hc25409e0} /* (8, 9, 10) {real, imag} */,
  {32'h42845f5d, 32'hc231de7f} /* (8, 9, 9) {real, imag} */,
  {32'h42c595b1, 32'hc1bb661e} /* (8, 9, 8) {real, imag} */,
  {32'hc26e9df5, 32'hc233ad71} /* (8, 9, 7) {real, imag} */,
  {32'h427db2c1, 32'hc1098261} /* (8, 9, 6) {real, imag} */,
  {32'hc32cc492, 32'hc2ae83ea} /* (8, 9, 5) {real, imag} */,
  {32'h43087d6a, 32'h42d388db} /* (8, 9, 4) {real, imag} */,
  {32'h4240d132, 32'h43125491} /* (8, 9, 3) {real, imag} */,
  {32'hc448360a, 32'hc3e03f2d} /* (8, 9, 2) {real, imag} */,
  {32'h44f30a1e, 32'h447e1134} /* (8, 9, 1) {real, imag} */,
  {32'h4506bc5c, 32'h00000000} /* (8, 9, 0) {real, imag} */,
  {32'h452d34cc, 32'hc4aca5d2} /* (8, 8, 31) {real, imag} */,
  {32'hc48695ba, 32'h4402ea10} /* (8, 8, 30) {real, imag} */,
  {32'h42d0de17, 32'hc22cec0f} /* (8, 8, 29) {real, imag} */,
  {32'h4300a73c, 32'hc2c220a0} /* (8, 8, 28) {real, imag} */,
  {32'hc320c182, 32'hc21ed40c} /* (8, 8, 27) {real, imag} */,
  {32'h42437d9e, 32'hc1cbaaf6} /* (8, 8, 26) {real, imag} */,
  {32'h418f8c10, 32'hc102431c} /* (8, 8, 25) {real, imag} */,
  {32'hc138b123, 32'h41e27e42} /* (8, 8, 24) {real, imag} */,
  {32'hc26aa5cc, 32'hc1da669c} /* (8, 8, 23) {real, imag} */,
  {32'h42a69046, 32'hc155ec56} /* (8, 8, 22) {real, imag} */,
  {32'h421f8678, 32'h41ec45be} /* (8, 8, 21) {real, imag} */,
  {32'h41d3645f, 32'hc24cea2a} /* (8, 8, 20) {real, imag} */,
  {32'hc296def2, 32'hc2553bec} /* (8, 8, 19) {real, imag} */,
  {32'hc3055c53, 32'hc1db169d} /* (8, 8, 18) {real, imag} */,
  {32'hc20f2ee8, 32'hc1974ffa} /* (8, 8, 17) {real, imag} */,
  {32'h42dfdead, 32'h00000000} /* (8, 8, 16) {real, imag} */,
  {32'hc20f2ee8, 32'h41974ffa} /* (8, 8, 15) {real, imag} */,
  {32'hc3055c53, 32'h41db169d} /* (8, 8, 14) {real, imag} */,
  {32'hc296def2, 32'h42553bec} /* (8, 8, 13) {real, imag} */,
  {32'h41d3645f, 32'h424cea2a} /* (8, 8, 12) {real, imag} */,
  {32'h421f8678, 32'hc1ec45be} /* (8, 8, 11) {real, imag} */,
  {32'h42a69046, 32'h4155ec56} /* (8, 8, 10) {real, imag} */,
  {32'hc26aa5cc, 32'h41da669c} /* (8, 8, 9) {real, imag} */,
  {32'hc138b123, 32'hc1e27e42} /* (8, 8, 8) {real, imag} */,
  {32'h418f8c10, 32'h4102431c} /* (8, 8, 7) {real, imag} */,
  {32'h42437d9e, 32'h41cbaaf6} /* (8, 8, 6) {real, imag} */,
  {32'hc320c182, 32'h421ed40c} /* (8, 8, 5) {real, imag} */,
  {32'h4300a73c, 32'h42c220a0} /* (8, 8, 4) {real, imag} */,
  {32'h42d0de17, 32'h422cec0f} /* (8, 8, 3) {real, imag} */,
  {32'hc48695ba, 32'hc402ea10} /* (8, 8, 2) {real, imag} */,
  {32'h452d34cc, 32'h44aca5d2} /* (8, 8, 1) {real, imag} */,
  {32'h4541489c, 32'h00000000} /* (8, 8, 0) {real, imag} */,
  {32'h454f2c10, 32'hc4ca0631} /* (8, 7, 31) {real, imag} */,
  {32'hc48e6964, 32'h4424ef50} /* (8, 7, 30) {real, imag} */,
  {32'h4303aa3f, 32'hc299b6c7} /* (8, 7, 29) {real, imag} */,
  {32'h43161424, 32'hc3019e10} /* (8, 7, 28) {real, imag} */,
  {32'hc383fd4a, 32'h432d89f1} /* (8, 7, 27) {real, imag} */,
  {32'hc2e68484, 32'h427e8cdf} /* (8, 7, 26) {real, imag} */,
  {32'h42c57f8a, 32'hc28890be} /* (8, 7, 25) {real, imag} */,
  {32'h429b7c12, 32'h42fca390} /* (8, 7, 24) {real, imag} */,
  {32'h420da715, 32'h4269acba} /* (8, 7, 23) {real, imag} */,
  {32'h41be6300, 32'h41bab8e4} /* (8, 7, 22) {real, imag} */,
  {32'h41e72e96, 32'h4209f32c} /* (8, 7, 21) {real, imag} */,
  {32'h42c3679e, 32'h41e61694} /* (8, 7, 20) {real, imag} */,
  {32'h42cbce5b, 32'hc22fa8bc} /* (8, 7, 19) {real, imag} */,
  {32'hc1bc1ed0, 32'h41f52536} /* (8, 7, 18) {real, imag} */,
  {32'hc29e2878, 32'hc261e02c} /* (8, 7, 17) {real, imag} */,
  {32'h419219c4, 32'h00000000} /* (8, 7, 16) {real, imag} */,
  {32'hc29e2878, 32'h4261e02c} /* (8, 7, 15) {real, imag} */,
  {32'hc1bc1ed0, 32'hc1f52536} /* (8, 7, 14) {real, imag} */,
  {32'h42cbce5b, 32'h422fa8bc} /* (8, 7, 13) {real, imag} */,
  {32'h42c3679e, 32'hc1e61694} /* (8, 7, 12) {real, imag} */,
  {32'h41e72e96, 32'hc209f32c} /* (8, 7, 11) {real, imag} */,
  {32'h41be6300, 32'hc1bab8e4} /* (8, 7, 10) {real, imag} */,
  {32'h420da715, 32'hc269acba} /* (8, 7, 9) {real, imag} */,
  {32'h429b7c12, 32'hc2fca390} /* (8, 7, 8) {real, imag} */,
  {32'h42c57f8a, 32'h428890be} /* (8, 7, 7) {real, imag} */,
  {32'hc2e68484, 32'hc27e8cdf} /* (8, 7, 6) {real, imag} */,
  {32'hc383fd4a, 32'hc32d89f1} /* (8, 7, 5) {real, imag} */,
  {32'h43161424, 32'h43019e10} /* (8, 7, 4) {real, imag} */,
  {32'h4303aa3f, 32'h4299b6c7} /* (8, 7, 3) {real, imag} */,
  {32'hc48e6964, 32'hc424ef50} /* (8, 7, 2) {real, imag} */,
  {32'h454f2c10, 32'h44ca0631} /* (8, 7, 1) {real, imag} */,
  {32'h456bc8bf, 32'h00000000} /* (8, 7, 0) {real, imag} */,
  {32'h455a8070, 32'hc5036202} /* (8, 6, 31) {real, imag} */,
  {32'hc46cddba, 32'h4459f31d} /* (8, 6, 30) {real, imag} */,
  {32'h40844aec, 32'hc1c25c5f} /* (8, 6, 29) {real, imag} */,
  {32'h42d8a4ec, 32'h4107c7a4} /* (8, 6, 28) {real, imag} */,
  {32'hc3586115, 32'h42efd4d4} /* (8, 6, 27) {real, imag} */,
  {32'h40d35428, 32'h422f071e} /* (8, 6, 26) {real, imag} */,
  {32'hc1a27d38, 32'hc241f7ce} /* (8, 6, 25) {real, imag} */,
  {32'hc29cac5a, 32'h424bb047} /* (8, 6, 24) {real, imag} */,
  {32'hc078288c, 32'hc234f296} /* (8, 6, 23) {real, imag} */,
  {32'hc281d17c, 32'hc201f455} /* (8, 6, 22) {real, imag} */,
  {32'h426cc484, 32'hc1e235ac} /* (8, 6, 21) {real, imag} */,
  {32'h415e70a8, 32'hc26a8daf} /* (8, 6, 20) {real, imag} */,
  {32'hc1a1e41b, 32'h419a6c05} /* (8, 6, 19) {real, imag} */,
  {32'hc0af089a, 32'hc1c7cb5e} /* (8, 6, 18) {real, imag} */,
  {32'h4275cffa, 32'hc1d8219d} /* (8, 6, 17) {real, imag} */,
  {32'h42be4cce, 32'h00000000} /* (8, 6, 16) {real, imag} */,
  {32'h4275cffa, 32'h41d8219d} /* (8, 6, 15) {real, imag} */,
  {32'hc0af089a, 32'h41c7cb5e} /* (8, 6, 14) {real, imag} */,
  {32'hc1a1e41b, 32'hc19a6c05} /* (8, 6, 13) {real, imag} */,
  {32'h415e70a8, 32'h426a8daf} /* (8, 6, 12) {real, imag} */,
  {32'h426cc484, 32'h41e235ac} /* (8, 6, 11) {real, imag} */,
  {32'hc281d17c, 32'h4201f455} /* (8, 6, 10) {real, imag} */,
  {32'hc078288c, 32'h4234f296} /* (8, 6, 9) {real, imag} */,
  {32'hc29cac5a, 32'hc24bb047} /* (8, 6, 8) {real, imag} */,
  {32'hc1a27d38, 32'h4241f7ce} /* (8, 6, 7) {real, imag} */,
  {32'h40d35428, 32'hc22f071e} /* (8, 6, 6) {real, imag} */,
  {32'hc3586115, 32'hc2efd4d4} /* (8, 6, 5) {real, imag} */,
  {32'h42d8a4ec, 32'hc107c7a4} /* (8, 6, 4) {real, imag} */,
  {32'h40844aec, 32'h41c25c5f} /* (8, 6, 3) {real, imag} */,
  {32'hc46cddba, 32'hc459f31d} /* (8, 6, 2) {real, imag} */,
  {32'h455a8070, 32'h45036202} /* (8, 6, 1) {real, imag} */,
  {32'h458310c7, 32'h00000000} /* (8, 6, 0) {real, imag} */,
  {32'h454e6375, 32'hc536f323} /* (8, 5, 31) {real, imag} */,
  {32'hc3c06df4, 32'h44868fe3} /* (8, 5, 30) {real, imag} */,
  {32'h427a81ed, 32'hc24a82ef} /* (8, 5, 29) {real, imag} */,
  {32'h3f721d00, 32'h43456a7a} /* (8, 5, 28) {real, imag} */,
  {32'hc26ff3a6, 32'h421114e8} /* (8, 5, 27) {real, imag} */,
  {32'h42b0765f, 32'h42c4a23a} /* (8, 5, 26) {real, imag} */,
  {32'h429679f0, 32'hc1478370} /* (8, 5, 25) {real, imag} */,
  {32'h429b35e2, 32'h42803424} /* (8, 5, 24) {real, imag} */,
  {32'h4113b33d, 32'h42f9cd01} /* (8, 5, 23) {real, imag} */,
  {32'h421e2012, 32'h42422c13} /* (8, 5, 22) {real, imag} */,
  {32'hc2c80992, 32'hc1e2755c} /* (8, 5, 21) {real, imag} */,
  {32'hc25ded4a, 32'hc20a5384} /* (8, 5, 20) {real, imag} */,
  {32'h42c047a7, 32'hc2b447d3} /* (8, 5, 19) {real, imag} */,
  {32'h41b50e9f, 32'h41187b41} /* (8, 5, 18) {real, imag} */,
  {32'hc2112556, 32'h42c6dcc5} /* (8, 5, 17) {real, imag} */,
  {32'hc2a9a751, 32'h00000000} /* (8, 5, 16) {real, imag} */,
  {32'hc2112556, 32'hc2c6dcc5} /* (8, 5, 15) {real, imag} */,
  {32'h41b50e9f, 32'hc1187b41} /* (8, 5, 14) {real, imag} */,
  {32'h42c047a7, 32'h42b447d3} /* (8, 5, 13) {real, imag} */,
  {32'hc25ded4a, 32'h420a5384} /* (8, 5, 12) {real, imag} */,
  {32'hc2c80992, 32'h41e2755c} /* (8, 5, 11) {real, imag} */,
  {32'h421e2012, 32'hc2422c13} /* (8, 5, 10) {real, imag} */,
  {32'h4113b33d, 32'hc2f9cd01} /* (8, 5, 9) {real, imag} */,
  {32'h429b35e2, 32'hc2803424} /* (8, 5, 8) {real, imag} */,
  {32'h429679f0, 32'h41478370} /* (8, 5, 7) {real, imag} */,
  {32'h42b0765f, 32'hc2c4a23a} /* (8, 5, 6) {real, imag} */,
  {32'hc26ff3a6, 32'hc21114e8} /* (8, 5, 5) {real, imag} */,
  {32'h3f721d00, 32'hc3456a7a} /* (8, 5, 4) {real, imag} */,
  {32'h427a81ed, 32'h424a82ef} /* (8, 5, 3) {real, imag} */,
  {32'hc3c06df4, 32'hc4868fe3} /* (8, 5, 2) {real, imag} */,
  {32'h454e6375, 32'h4536f323} /* (8, 5, 1) {real, imag} */,
  {32'h4599ba1a, 32'h00000000} /* (8, 5, 0) {real, imag} */,
  {32'h453bcf36, 32'hc54f89b0} /* (8, 4, 31) {real, imag} */,
  {32'h424a4ff0, 32'h4493e68e} /* (8, 4, 30) {real, imag} */,
  {32'hc244aa1c, 32'h422c56cb} /* (8, 4, 29) {real, imag} */,
  {32'hc2c6b56c, 32'h434dcf19} /* (8, 4, 28) {real, imag} */,
  {32'hc3044de0, 32'h42c42dc3} /* (8, 4, 27) {real, imag} */,
  {32'h42a22480, 32'h42ab28a2} /* (8, 4, 26) {real, imag} */,
  {32'h4298dba4, 32'hc2e59b20} /* (8, 4, 25) {real, imag} */,
  {32'hc085c380, 32'h420438cb} /* (8, 4, 24) {real, imag} */,
  {32'hc231a829, 32'hc2eae782} /* (8, 4, 23) {real, imag} */,
  {32'hc1e8163a, 32'h42c53832} /* (8, 4, 22) {real, imag} */,
  {32'hc305124d, 32'h41938314} /* (8, 4, 21) {real, imag} */,
  {32'h422812bd, 32'h4259e0e4} /* (8, 4, 20) {real, imag} */,
  {32'h428e14e5, 32'h41d3e8e4} /* (8, 4, 19) {real, imag} */,
  {32'h420b8b30, 32'h400ae638} /* (8, 4, 18) {real, imag} */,
  {32'hc24235cf, 32'h41e12ee8} /* (8, 4, 17) {real, imag} */,
  {32'hbdeb3c00, 32'h00000000} /* (8, 4, 16) {real, imag} */,
  {32'hc24235cf, 32'hc1e12ee8} /* (8, 4, 15) {real, imag} */,
  {32'h420b8b30, 32'hc00ae638} /* (8, 4, 14) {real, imag} */,
  {32'h428e14e5, 32'hc1d3e8e4} /* (8, 4, 13) {real, imag} */,
  {32'h422812bd, 32'hc259e0e4} /* (8, 4, 12) {real, imag} */,
  {32'hc305124d, 32'hc1938314} /* (8, 4, 11) {real, imag} */,
  {32'hc1e8163a, 32'hc2c53832} /* (8, 4, 10) {real, imag} */,
  {32'hc231a829, 32'h42eae782} /* (8, 4, 9) {real, imag} */,
  {32'hc085c380, 32'hc20438cb} /* (8, 4, 8) {real, imag} */,
  {32'h4298dba4, 32'h42e59b20} /* (8, 4, 7) {real, imag} */,
  {32'h42a22480, 32'hc2ab28a2} /* (8, 4, 6) {real, imag} */,
  {32'hc3044de0, 32'hc2c42dc3} /* (8, 4, 5) {real, imag} */,
  {32'hc2c6b56c, 32'hc34dcf19} /* (8, 4, 4) {real, imag} */,
  {32'hc244aa1c, 32'hc22c56cb} /* (8, 4, 3) {real, imag} */,
  {32'h424a4ff0, 32'hc493e68e} /* (8, 4, 2) {real, imag} */,
  {32'h453bcf36, 32'h454f89b0} /* (8, 4, 1) {real, imag} */,
  {32'h45a36678, 32'h00000000} /* (8, 4, 0) {real, imag} */,
  {32'h45376d5e, 32'hc563b414} /* (8, 3, 31) {real, imag} */,
  {32'h4372fcb0, 32'h44898a86} /* (8, 3, 30) {real, imag} */,
  {32'hc2930fd8, 32'h42c6ccb0} /* (8, 3, 29) {real, imag} */,
  {32'hc2379860, 32'h439e024e} /* (8, 3, 28) {real, imag} */,
  {32'hc31a1852, 32'hc26c987e} /* (8, 3, 27) {real, imag} */,
  {32'hc2a6b8dc, 32'hc321c094} /* (8, 3, 26) {real, imag} */,
  {32'h41b0a260, 32'h42781dd6} /* (8, 3, 25) {real, imag} */,
  {32'hc1dc41a4, 32'h41d020f7} /* (8, 3, 24) {real, imag} */,
  {32'h42cb902c, 32'h41c86c4c} /* (8, 3, 23) {real, imag} */,
  {32'hc262d00c, 32'h42b6c78c} /* (8, 3, 22) {real, imag} */,
  {32'hc27f660d, 32'hbfc06680} /* (8, 3, 21) {real, imag} */,
  {32'h43102309, 32'h40b834fa} /* (8, 3, 20) {real, imag} */,
  {32'hc2b2b26f, 32'h40c16870} /* (8, 3, 19) {real, imag} */,
  {32'hc24daa98, 32'h4204e9f5} /* (8, 3, 18) {real, imag} */,
  {32'hc1e0302c, 32'h4141bb44} /* (8, 3, 17) {real, imag} */,
  {32'hc2966662, 32'h00000000} /* (8, 3, 16) {real, imag} */,
  {32'hc1e0302c, 32'hc141bb44} /* (8, 3, 15) {real, imag} */,
  {32'hc24daa98, 32'hc204e9f5} /* (8, 3, 14) {real, imag} */,
  {32'hc2b2b26f, 32'hc0c16870} /* (8, 3, 13) {real, imag} */,
  {32'h43102309, 32'hc0b834fa} /* (8, 3, 12) {real, imag} */,
  {32'hc27f660d, 32'h3fc06680} /* (8, 3, 11) {real, imag} */,
  {32'hc262d00c, 32'hc2b6c78c} /* (8, 3, 10) {real, imag} */,
  {32'h42cb902c, 32'hc1c86c4c} /* (8, 3, 9) {real, imag} */,
  {32'hc1dc41a4, 32'hc1d020f7} /* (8, 3, 8) {real, imag} */,
  {32'h41b0a260, 32'hc2781dd6} /* (8, 3, 7) {real, imag} */,
  {32'hc2a6b8dc, 32'h4321c094} /* (8, 3, 6) {real, imag} */,
  {32'hc31a1852, 32'h426c987e} /* (8, 3, 5) {real, imag} */,
  {32'hc2379860, 32'hc39e024e} /* (8, 3, 4) {real, imag} */,
  {32'hc2930fd8, 32'hc2c6ccb0} /* (8, 3, 3) {real, imag} */,
  {32'h4372fcb0, 32'hc4898a86} /* (8, 3, 2) {real, imag} */,
  {32'h45376d5e, 32'h4563b414} /* (8, 3, 1) {real, imag} */,
  {32'h45a4409b, 32'h00000000} /* (8, 3, 0) {real, imag} */,
  {32'h453c7398, 32'hc566e3be} /* (8, 2, 31) {real, imag} */,
  {32'h43d12c91, 32'h44904aaa} /* (8, 2, 30) {real, imag} */,
  {32'hc3524b9b, 32'h4383b49d} /* (8, 2, 29) {real, imag} */,
  {32'hc2ca7ed7, 32'h438cfafb} /* (8, 2, 28) {real, imag} */,
  {32'hc3207806, 32'hc3317201} /* (8, 2, 27) {real, imag} */,
  {32'hc230fabc, 32'hc199d881} /* (8, 2, 26) {real, imag} */,
  {32'h40fcd010, 32'h4258de1d} /* (8, 2, 25) {real, imag} */,
  {32'h42df1424, 32'h41ff4c00} /* (8, 2, 24) {real, imag} */,
  {32'hc279b024, 32'h430fc2f4} /* (8, 2, 23) {real, imag} */,
  {32'hc28f6b3e, 32'h42ced0cd} /* (8, 2, 22) {real, imag} */,
  {32'hc2bd0b64, 32'hc2d47202} /* (8, 2, 21) {real, imag} */,
  {32'h4128d906, 32'hc28bea5e} /* (8, 2, 20) {real, imag} */,
  {32'h421a0d26, 32'hc28fe42c} /* (8, 2, 19) {real, imag} */,
  {32'h41ad108f, 32'h42dbd03e} /* (8, 2, 18) {real, imag} */,
  {32'hc114b2bf, 32'h423d1a2e} /* (8, 2, 17) {real, imag} */,
  {32'hc29ec37e, 32'h00000000} /* (8, 2, 16) {real, imag} */,
  {32'hc114b2bf, 32'hc23d1a2e} /* (8, 2, 15) {real, imag} */,
  {32'h41ad108f, 32'hc2dbd03e} /* (8, 2, 14) {real, imag} */,
  {32'h421a0d26, 32'h428fe42c} /* (8, 2, 13) {real, imag} */,
  {32'h4128d906, 32'h428bea5e} /* (8, 2, 12) {real, imag} */,
  {32'hc2bd0b64, 32'h42d47202} /* (8, 2, 11) {real, imag} */,
  {32'hc28f6b3e, 32'hc2ced0cd} /* (8, 2, 10) {real, imag} */,
  {32'hc279b024, 32'hc30fc2f4} /* (8, 2, 9) {real, imag} */,
  {32'h42df1424, 32'hc1ff4c00} /* (8, 2, 8) {real, imag} */,
  {32'h40fcd010, 32'hc258de1d} /* (8, 2, 7) {real, imag} */,
  {32'hc230fabc, 32'h4199d881} /* (8, 2, 6) {real, imag} */,
  {32'hc3207806, 32'h43317201} /* (8, 2, 5) {real, imag} */,
  {32'hc2ca7ed7, 32'hc38cfafb} /* (8, 2, 4) {real, imag} */,
  {32'hc3524b9b, 32'hc383b49d} /* (8, 2, 3) {real, imag} */,
  {32'h43d12c91, 32'hc4904aaa} /* (8, 2, 2) {real, imag} */,
  {32'h453c7398, 32'h4566e3be} /* (8, 2, 1) {real, imag} */,
  {32'h45aa85c8, 32'h00000000} /* (8, 2, 0) {real, imag} */,
  {32'h453e08cb, 32'hc553afb8} /* (8, 1, 31) {real, imag} */,
  {32'h43555dd2, 32'h446477b2} /* (8, 1, 30) {real, imag} */,
  {32'hc3767c2c, 32'h4346b20d} /* (8, 1, 29) {real, imag} */,
  {32'hc26b0f6b, 32'h43a55397} /* (8, 1, 28) {real, imag} */,
  {32'hc2ca4b50, 32'hc2f60fc3} /* (8, 1, 27) {real, imag} */,
  {32'h4041ac28, 32'hc235718a} /* (8, 1, 26) {real, imag} */,
  {32'hc2a4cb13, 32'h42844bea} /* (8, 1, 25) {real, imag} */,
  {32'h42a07628, 32'hc1e3e90b} /* (8, 1, 24) {real, imag} */,
  {32'hc12ca7a2, 32'hc215d356} /* (8, 1, 23) {real, imag} */,
  {32'h407a3a40, 32'h42b809a4} /* (8, 1, 22) {real, imag} */,
  {32'hc280baea, 32'hbfb5ce20} /* (8, 1, 21) {real, imag} */,
  {32'h42a1bb28, 32'hc2d3f0b1} /* (8, 1, 20) {real, imag} */,
  {32'h41bbb750, 32'h42b21b4e} /* (8, 1, 19) {real, imag} */,
  {32'hc110fc1c, 32'hc19248a6} /* (8, 1, 18) {real, imag} */,
  {32'hc1a7f013, 32'hc205877a} /* (8, 1, 17) {real, imag} */,
  {32'hc1ac4d0a, 32'h00000000} /* (8, 1, 16) {real, imag} */,
  {32'hc1a7f013, 32'h4205877a} /* (8, 1, 15) {real, imag} */,
  {32'hc110fc1c, 32'h419248a6} /* (8, 1, 14) {real, imag} */,
  {32'h41bbb750, 32'hc2b21b4e} /* (8, 1, 13) {real, imag} */,
  {32'h42a1bb28, 32'h42d3f0b1} /* (8, 1, 12) {real, imag} */,
  {32'hc280baea, 32'h3fb5ce20} /* (8, 1, 11) {real, imag} */,
  {32'h407a3a40, 32'hc2b809a4} /* (8, 1, 10) {real, imag} */,
  {32'hc12ca7a2, 32'h4215d356} /* (8, 1, 9) {real, imag} */,
  {32'h42a07628, 32'h41e3e90b} /* (8, 1, 8) {real, imag} */,
  {32'hc2a4cb13, 32'hc2844bea} /* (8, 1, 7) {real, imag} */,
  {32'h4041ac28, 32'h4235718a} /* (8, 1, 6) {real, imag} */,
  {32'hc2ca4b50, 32'h42f60fc3} /* (8, 1, 5) {real, imag} */,
  {32'hc26b0f6b, 32'hc3a55397} /* (8, 1, 4) {real, imag} */,
  {32'hc3767c2c, 32'hc346b20d} /* (8, 1, 3) {real, imag} */,
  {32'h43555dd2, 32'hc46477b2} /* (8, 1, 2) {real, imag} */,
  {32'h453e08cb, 32'h4553afb8} /* (8, 1, 1) {real, imag} */,
  {32'h45a7271f, 32'h00000000} /* (8, 1, 0) {real, imag} */,
  {32'h454677d7, 32'hc52ede9a} /* (8, 0, 31) {real, imag} */,
  {32'hc2a4bcc8, 32'h443c6c82} /* (8, 0, 30) {real, imag} */,
  {32'hc35dafcc, 32'h42b2c60e} /* (8, 0, 29) {real, imag} */,
  {32'h40ebb548, 32'h4377fc34} /* (8, 0, 28) {real, imag} */,
  {32'hc2a01cdc, 32'hc2d6c1f9} /* (8, 0, 27) {real, imag} */,
  {32'hc1fde1b8, 32'h4208944c} /* (8, 0, 26) {real, imag} */,
  {32'hc2845720, 32'hbef4f340} /* (8, 0, 25) {real, imag} */,
  {32'h41904328, 32'h4185d1ce} /* (8, 0, 24) {real, imag} */,
  {32'h3caa2800, 32'h4146b4c0} /* (8, 0, 23) {real, imag} */,
  {32'hc1bfd260, 32'hc22b460f} /* (8, 0, 22) {real, imag} */,
  {32'h421bd0ff, 32'h428d58b7} /* (8, 0, 21) {real, imag} */,
  {32'h42f23c2e, 32'h40cc47c0} /* (8, 0, 20) {real, imag} */,
  {32'hbdda0d00, 32'hc1a4a8a2} /* (8, 0, 19) {real, imag} */,
  {32'hc20a9f6b, 32'hc2420cbc} /* (8, 0, 18) {real, imag} */,
  {32'h4181a0e6, 32'h424038b4} /* (8, 0, 17) {real, imag} */,
  {32'hc24c8d7d, 32'h00000000} /* (8, 0, 16) {real, imag} */,
  {32'h4181a0e6, 32'hc24038b4} /* (8, 0, 15) {real, imag} */,
  {32'hc20a9f6b, 32'h42420cbc} /* (8, 0, 14) {real, imag} */,
  {32'hbdda0d00, 32'h41a4a8a2} /* (8, 0, 13) {real, imag} */,
  {32'h42f23c2e, 32'hc0cc47c0} /* (8, 0, 12) {real, imag} */,
  {32'h421bd0ff, 32'hc28d58b7} /* (8, 0, 11) {real, imag} */,
  {32'hc1bfd260, 32'h422b460f} /* (8, 0, 10) {real, imag} */,
  {32'h3caa2800, 32'hc146b4c0} /* (8, 0, 9) {real, imag} */,
  {32'h41904328, 32'hc185d1ce} /* (8, 0, 8) {real, imag} */,
  {32'hc2845720, 32'h3ef4f340} /* (8, 0, 7) {real, imag} */,
  {32'hc1fde1b8, 32'hc208944c} /* (8, 0, 6) {real, imag} */,
  {32'hc2a01cdc, 32'h42d6c1f9} /* (8, 0, 5) {real, imag} */,
  {32'h40ebb548, 32'hc377fc34} /* (8, 0, 4) {real, imag} */,
  {32'hc35dafcc, 32'hc2b2c60e} /* (8, 0, 3) {real, imag} */,
  {32'hc2a4bcc8, 32'hc43c6c82} /* (8, 0, 2) {real, imag} */,
  {32'h454677d7, 32'h452ede9a} /* (8, 0, 1) {real, imag} */,
  {32'h45a025b5, 32'h00000000} /* (8, 0, 0) {real, imag} */,
  {32'h4540025a, 32'hc4ccfbe4} /* (7, 31, 31) {real, imag} */,
  {32'hc3ec3489, 32'h43c0bdeb} /* (7, 31, 30) {real, imag} */,
  {32'hc2b4f2fb, 32'h40eaf3d0} /* (7, 31, 29) {real, imag} */,
  {32'h4312c268, 32'h41eb6df0} /* (7, 31, 28) {real, imag} */,
  {32'hc2db0233, 32'h42377c51} /* (7, 31, 27) {real, imag} */,
  {32'h402d1100, 32'h42168f05} /* (7, 31, 26) {real, imag} */,
  {32'h4117efad, 32'h4237c9c9} /* (7, 31, 25) {real, imag} */,
  {32'hc2e83951, 32'h422a9963} /* (7, 31, 24) {real, imag} */,
  {32'h4263eb56, 32'hc235ff9b} /* (7, 31, 23) {real, imag} */,
  {32'h42a164a9, 32'h429577e8} /* (7, 31, 22) {real, imag} */,
  {32'hc2b53de8, 32'h428863c6} /* (7, 31, 21) {real, imag} */,
  {32'hc1e2382a, 32'hc21800f8} /* (7, 31, 20) {real, imag} */,
  {32'h41975308, 32'hc18544ab} /* (7, 31, 19) {real, imag} */,
  {32'h41d69e92, 32'h424437a9} /* (7, 31, 18) {real, imag} */,
  {32'hc1c38a32, 32'h419082b2} /* (7, 31, 17) {real, imag} */,
  {32'hc2b7ead1, 32'h00000000} /* (7, 31, 16) {real, imag} */,
  {32'hc1c38a32, 32'hc19082b2} /* (7, 31, 15) {real, imag} */,
  {32'h41d69e92, 32'hc24437a9} /* (7, 31, 14) {real, imag} */,
  {32'h41975308, 32'h418544ab} /* (7, 31, 13) {real, imag} */,
  {32'hc1e2382a, 32'h421800f8} /* (7, 31, 12) {real, imag} */,
  {32'hc2b53de8, 32'hc28863c6} /* (7, 31, 11) {real, imag} */,
  {32'h42a164a9, 32'hc29577e8} /* (7, 31, 10) {real, imag} */,
  {32'h4263eb56, 32'h4235ff9b} /* (7, 31, 9) {real, imag} */,
  {32'hc2e83951, 32'hc22a9963} /* (7, 31, 8) {real, imag} */,
  {32'h4117efad, 32'hc237c9c9} /* (7, 31, 7) {real, imag} */,
  {32'h402d1100, 32'hc2168f05} /* (7, 31, 6) {real, imag} */,
  {32'hc2db0233, 32'hc2377c51} /* (7, 31, 5) {real, imag} */,
  {32'h4312c268, 32'hc1eb6df0} /* (7, 31, 4) {real, imag} */,
  {32'hc2b4f2fb, 32'hc0eaf3d0} /* (7, 31, 3) {real, imag} */,
  {32'hc3ec3489, 32'hc3c0bdeb} /* (7, 31, 2) {real, imag} */,
  {32'h4540025a, 32'h44ccfbe4} /* (7, 31, 1) {real, imag} */,
  {32'h458c1258, 32'h00000000} /* (7, 31, 0) {real, imag} */,
  {32'h4566b534, 32'hc49a89d2} /* (7, 30, 31) {real, imag} */,
  {32'hc455c914, 32'h43d71557} /* (7, 30, 30) {real, imag} */,
  {32'hc1e77864, 32'h42aaa002} /* (7, 30, 29) {real, imag} */,
  {32'h4324195a, 32'hc3012400} /* (7, 30, 28) {real, imag} */,
  {32'hc384f0dd, 32'h42a43f2e} /* (7, 30, 27) {real, imag} */,
  {32'hc228bcbf, 32'h432ace48} /* (7, 30, 26) {real, imag} */,
  {32'h42c944b6, 32'hc1b6d44a} /* (7, 30, 25) {real, imag} */,
  {32'hc2f09a0e, 32'h424c3864} /* (7, 30, 24) {real, imag} */,
  {32'hbf8171e0, 32'h42833542} /* (7, 30, 23) {real, imag} */,
  {32'hc13646ea, 32'hc0eb80a8} /* (7, 30, 22) {real, imag} */,
  {32'hc2a241c0, 32'h40689c40} /* (7, 30, 21) {real, imag} */,
  {32'hc2748f62, 32'hc20c0e6c} /* (7, 30, 20) {real, imag} */,
  {32'hc138de26, 32'hc1986310} /* (7, 30, 19) {real, imag} */,
  {32'hc21c8da4, 32'hc1eaddf0} /* (7, 30, 18) {real, imag} */,
  {32'h426a5251, 32'hc2c1e4b8} /* (7, 30, 17) {real, imag} */,
  {32'h41465dce, 32'h00000000} /* (7, 30, 16) {real, imag} */,
  {32'h426a5251, 32'h42c1e4b8} /* (7, 30, 15) {real, imag} */,
  {32'hc21c8da4, 32'h41eaddf0} /* (7, 30, 14) {real, imag} */,
  {32'hc138de26, 32'h41986310} /* (7, 30, 13) {real, imag} */,
  {32'hc2748f62, 32'h420c0e6c} /* (7, 30, 12) {real, imag} */,
  {32'hc2a241c0, 32'hc0689c40} /* (7, 30, 11) {real, imag} */,
  {32'hc13646ea, 32'h40eb80a8} /* (7, 30, 10) {real, imag} */,
  {32'hbf8171e0, 32'hc2833542} /* (7, 30, 9) {real, imag} */,
  {32'hc2f09a0e, 32'hc24c3864} /* (7, 30, 8) {real, imag} */,
  {32'h42c944b6, 32'h41b6d44a} /* (7, 30, 7) {real, imag} */,
  {32'hc228bcbf, 32'hc32ace48} /* (7, 30, 6) {real, imag} */,
  {32'hc384f0dd, 32'hc2a43f2e} /* (7, 30, 5) {real, imag} */,
  {32'h4324195a, 32'h43012400} /* (7, 30, 4) {real, imag} */,
  {32'hc1e77864, 32'hc2aaa002} /* (7, 30, 3) {real, imag} */,
  {32'hc455c914, 32'hc3d71557} /* (7, 30, 2) {real, imag} */,
  {32'h4566b534, 32'h449a89d2} /* (7, 30, 1) {real, imag} */,
  {32'h458b44fc, 32'h00000000} /* (7, 30, 0) {real, imag} */,
  {32'h4572cff6, 32'hc440404c} /* (7, 29, 31) {real, imag} */,
  {32'hc477c517, 32'h43eae323} /* (7, 29, 30) {real, imag} */,
  {32'hc2511e34, 32'h42645fce} /* (7, 29, 29) {real, imag} */,
  {32'h4325b38e, 32'hc189ccf8} /* (7, 29, 28) {real, imag} */,
  {32'hc387f5f2, 32'h4298ad13} /* (7, 29, 27) {real, imag} */,
  {32'h4187c220, 32'h4248adfe} /* (7, 29, 26) {real, imag} */,
  {32'h424804fc, 32'hc2a3b22e} /* (7, 29, 25) {real, imag} */,
  {32'hc2d521b9, 32'h430b633c} /* (7, 29, 24) {real, imag} */,
  {32'h4192e01a, 32'h41d09525} /* (7, 29, 23) {real, imag} */,
  {32'hc1fefcc0, 32'hc2f88288} /* (7, 29, 22) {real, imag} */,
  {32'hc21fa45a, 32'h420b30a7} /* (7, 29, 21) {real, imag} */,
  {32'h42cb71f2, 32'hc25d91c4} /* (7, 29, 20) {real, imag} */,
  {32'hc1b90438, 32'hc0e1c160} /* (7, 29, 19) {real, imag} */,
  {32'h422acae6, 32'h42b169dc} /* (7, 29, 18) {real, imag} */,
  {32'h42384e3f, 32'hc284bdd8} /* (7, 29, 17) {real, imag} */,
  {32'hc1f75012, 32'h00000000} /* (7, 29, 16) {real, imag} */,
  {32'h42384e3f, 32'h4284bdd8} /* (7, 29, 15) {real, imag} */,
  {32'h422acae6, 32'hc2b169dc} /* (7, 29, 14) {real, imag} */,
  {32'hc1b90438, 32'h40e1c160} /* (7, 29, 13) {real, imag} */,
  {32'h42cb71f2, 32'h425d91c4} /* (7, 29, 12) {real, imag} */,
  {32'hc21fa45a, 32'hc20b30a7} /* (7, 29, 11) {real, imag} */,
  {32'hc1fefcc0, 32'h42f88288} /* (7, 29, 10) {real, imag} */,
  {32'h4192e01a, 32'hc1d09525} /* (7, 29, 9) {real, imag} */,
  {32'hc2d521b9, 32'hc30b633c} /* (7, 29, 8) {real, imag} */,
  {32'h424804fc, 32'h42a3b22e} /* (7, 29, 7) {real, imag} */,
  {32'h4187c220, 32'hc248adfe} /* (7, 29, 6) {real, imag} */,
  {32'hc387f5f2, 32'hc298ad13} /* (7, 29, 5) {real, imag} */,
  {32'h4325b38e, 32'h4189ccf8} /* (7, 29, 4) {real, imag} */,
  {32'hc2511e34, 32'hc2645fce} /* (7, 29, 3) {real, imag} */,
  {32'hc477c517, 32'hc3eae323} /* (7, 29, 2) {real, imag} */,
  {32'h4572cff6, 32'h4440404c} /* (7, 29, 1) {real, imag} */,
  {32'h458b4dfb, 32'h00000000} /* (7, 29, 0) {real, imag} */,
  {32'h4568e901, 32'hc427cc3c} /* (7, 28, 31) {real, imag} */,
  {32'hc487abe7, 32'h43d434c7} /* (7, 28, 30) {real, imag} */,
  {32'hc1e5e9b0, 32'hc2ac738f} /* (7, 28, 29) {real, imag} */,
  {32'h429a17c3, 32'hc2f52f09} /* (7, 28, 28) {real, imag} */,
  {32'hc3473112, 32'h4261971a} /* (7, 28, 27) {real, imag} */,
  {32'hc255064d, 32'h41eab5f4} /* (7, 28, 26) {real, imag} */,
  {32'hc2338e4c, 32'hc0f79f20} /* (7, 28, 25) {real, imag} */,
  {32'h4293d0be, 32'hc144ab5e} /* (7, 28, 24) {real, imag} */,
  {32'h42188fc4, 32'hc1ca0def} /* (7, 28, 23) {real, imag} */,
  {32'h429e6f4e, 32'hc25dbb3e} /* (7, 28, 22) {real, imag} */,
  {32'hc2127367, 32'hc1362100} /* (7, 28, 21) {real, imag} */,
  {32'hc2452726, 32'hc1d67d66} /* (7, 28, 20) {real, imag} */,
  {32'hc2307b57, 32'hc25909e5} /* (7, 28, 19) {real, imag} */,
  {32'h42966db5, 32'h428151f0} /* (7, 28, 18) {real, imag} */,
  {32'hc1885d8c, 32'h42c529dc} /* (7, 28, 17) {real, imag} */,
  {32'hc232e5bc, 32'h00000000} /* (7, 28, 16) {real, imag} */,
  {32'hc1885d8c, 32'hc2c529dc} /* (7, 28, 15) {real, imag} */,
  {32'h42966db5, 32'hc28151f0} /* (7, 28, 14) {real, imag} */,
  {32'hc2307b57, 32'h425909e5} /* (7, 28, 13) {real, imag} */,
  {32'hc2452726, 32'h41d67d66} /* (7, 28, 12) {real, imag} */,
  {32'hc2127367, 32'h41362100} /* (7, 28, 11) {real, imag} */,
  {32'h429e6f4e, 32'h425dbb3e} /* (7, 28, 10) {real, imag} */,
  {32'h42188fc4, 32'h41ca0def} /* (7, 28, 9) {real, imag} */,
  {32'h4293d0be, 32'h4144ab5e} /* (7, 28, 8) {real, imag} */,
  {32'hc2338e4c, 32'h40f79f20} /* (7, 28, 7) {real, imag} */,
  {32'hc255064d, 32'hc1eab5f4} /* (7, 28, 6) {real, imag} */,
  {32'hc3473112, 32'hc261971a} /* (7, 28, 5) {real, imag} */,
  {32'h429a17c3, 32'h42f52f09} /* (7, 28, 4) {real, imag} */,
  {32'hc1e5e9b0, 32'h42ac738f} /* (7, 28, 3) {real, imag} */,
  {32'hc487abe7, 32'hc3d434c7} /* (7, 28, 2) {real, imag} */,
  {32'h4568e901, 32'h4427cc3c} /* (7, 28, 1) {real, imag} */,
  {32'h458b3e54, 32'h00000000} /* (7, 28, 0) {real, imag} */,
  {32'h456b4ea4, 32'hc4181e02} /* (7, 27, 31) {real, imag} */,
  {32'hc49be5a2, 32'h43bbb596} /* (7, 27, 30) {real, imag} */,
  {32'hc0d8bfbc, 32'hc1e5ec5d} /* (7, 27, 29) {real, imag} */,
  {32'h432cf618, 32'hc30d2dca} /* (7, 27, 28) {real, imag} */,
  {32'hc341356e, 32'h428900da} /* (7, 27, 27) {real, imag} */,
  {32'hc20e69cb, 32'hc1b0c138} /* (7, 27, 26) {real, imag} */,
  {32'h43080b78, 32'hc28e0415} /* (7, 27, 25) {real, imag} */,
  {32'h3dd1e200, 32'hc08b5bb0} /* (7, 27, 24) {real, imag} */,
  {32'h41adebfa, 32'hc2525cdc} /* (7, 27, 23) {real, imag} */,
  {32'hc114885e, 32'hc11fe0ae} /* (7, 27, 22) {real, imag} */,
  {32'hc1f08534, 32'h429b34b4} /* (7, 27, 21) {real, imag} */,
  {32'hc1591ec2, 32'hc280e4ed} /* (7, 27, 20) {real, imag} */,
  {32'hc1f26f8e, 32'hc2918150} /* (7, 27, 19) {real, imag} */,
  {32'hc1ecbb64, 32'h42a83bce} /* (7, 27, 18) {real, imag} */,
  {32'hc089822c, 32'h4217f8f1} /* (7, 27, 17) {real, imag} */,
  {32'hc1512d1a, 32'h00000000} /* (7, 27, 16) {real, imag} */,
  {32'hc089822c, 32'hc217f8f1} /* (7, 27, 15) {real, imag} */,
  {32'hc1ecbb64, 32'hc2a83bce} /* (7, 27, 14) {real, imag} */,
  {32'hc1f26f8e, 32'h42918150} /* (7, 27, 13) {real, imag} */,
  {32'hc1591ec2, 32'h4280e4ed} /* (7, 27, 12) {real, imag} */,
  {32'hc1f08534, 32'hc29b34b4} /* (7, 27, 11) {real, imag} */,
  {32'hc114885e, 32'h411fe0ae} /* (7, 27, 10) {real, imag} */,
  {32'h41adebfa, 32'h42525cdc} /* (7, 27, 9) {real, imag} */,
  {32'h3dd1e200, 32'h408b5bb0} /* (7, 27, 8) {real, imag} */,
  {32'h43080b78, 32'h428e0415} /* (7, 27, 7) {real, imag} */,
  {32'hc20e69cb, 32'h41b0c138} /* (7, 27, 6) {real, imag} */,
  {32'hc341356e, 32'hc28900da} /* (7, 27, 5) {real, imag} */,
  {32'h432cf618, 32'h430d2dca} /* (7, 27, 4) {real, imag} */,
  {32'hc0d8bfbc, 32'h41e5ec5d} /* (7, 27, 3) {real, imag} */,
  {32'hc49be5a2, 32'hc3bbb596} /* (7, 27, 2) {real, imag} */,
  {32'h456b4ea4, 32'h44181e02} /* (7, 27, 1) {real, imag} */,
  {32'h4584142f, 32'h00000000} /* (7, 27, 0) {real, imag} */,
  {32'h45635b62, 32'hc41e0339} /* (7, 26, 31) {real, imag} */,
  {32'hc4a7e94e, 32'h4362ae04} /* (7, 26, 30) {real, imag} */,
  {32'h42855c09, 32'hc2a3a92e} /* (7, 26, 29) {real, imag} */,
  {32'h42ddb3c7, 32'h4240f13b} /* (7, 26, 28) {real, imag} */,
  {32'hc33f86f9, 32'h427ab970} /* (7, 26, 27) {real, imag} */,
  {32'h4247156c, 32'h411a5070} /* (7, 26, 26) {real, imag} */,
  {32'h42b71dfb, 32'hc1e55240} /* (7, 26, 25) {real, imag} */,
  {32'h41904280, 32'h42c8635a} /* (7, 26, 24) {real, imag} */,
  {32'h42edfa52, 32'h42311cbf} /* (7, 26, 23) {real, imag} */,
  {32'h40949020, 32'hc1c7f18c} /* (7, 26, 22) {real, imag} */,
  {32'h4290585e, 32'h42542a37} /* (7, 26, 21) {real, imag} */,
  {32'h40d19c18, 32'h4111f58a} /* (7, 26, 20) {real, imag} */,
  {32'h4225fe36, 32'hc18472c1} /* (7, 26, 19) {real, imag} */,
  {32'h41191008, 32'h41767270} /* (7, 26, 18) {real, imag} */,
  {32'h41481f9a, 32'h416ab9c8} /* (7, 26, 17) {real, imag} */,
  {32'hc2761b5a, 32'h00000000} /* (7, 26, 16) {real, imag} */,
  {32'h41481f9a, 32'hc16ab9c8} /* (7, 26, 15) {real, imag} */,
  {32'h41191008, 32'hc1767270} /* (7, 26, 14) {real, imag} */,
  {32'h4225fe36, 32'h418472c1} /* (7, 26, 13) {real, imag} */,
  {32'h40d19c18, 32'hc111f58a} /* (7, 26, 12) {real, imag} */,
  {32'h4290585e, 32'hc2542a37} /* (7, 26, 11) {real, imag} */,
  {32'h40949020, 32'h41c7f18c} /* (7, 26, 10) {real, imag} */,
  {32'h42edfa52, 32'hc2311cbf} /* (7, 26, 9) {real, imag} */,
  {32'h41904280, 32'hc2c8635a} /* (7, 26, 8) {real, imag} */,
  {32'h42b71dfb, 32'h41e55240} /* (7, 26, 7) {real, imag} */,
  {32'h4247156c, 32'hc11a5070} /* (7, 26, 6) {real, imag} */,
  {32'hc33f86f9, 32'hc27ab970} /* (7, 26, 5) {real, imag} */,
  {32'h42ddb3c7, 32'hc240f13b} /* (7, 26, 4) {real, imag} */,
  {32'h42855c09, 32'h42a3a92e} /* (7, 26, 3) {real, imag} */,
  {32'hc4a7e94e, 32'hc362ae04} /* (7, 26, 2) {real, imag} */,
  {32'h45635b62, 32'h441e0339} /* (7, 26, 1) {real, imag} */,
  {32'h457ea796, 32'h00000000} /* (7, 26, 0) {real, imag} */,
  {32'h4552f8ef, 32'hc40d4b01} /* (7, 25, 31) {real, imag} */,
  {32'hc4aa006c, 32'h43532284} /* (7, 25, 30) {real, imag} */,
  {32'hc1b37b88, 32'hc2f19597} /* (7, 25, 29) {real, imag} */,
  {32'h4341f538, 32'hc17e0be8} /* (7, 25, 28) {real, imag} */,
  {32'hc34a75f3, 32'h42e9cf4c} /* (7, 25, 27) {real, imag} */,
  {32'h41b92754, 32'hc1b49783} /* (7, 25, 26) {real, imag} */,
  {32'h416a8085, 32'hc30f02cc} /* (7, 25, 25) {real, imag} */,
  {32'hc187c573, 32'h4216c24f} /* (7, 25, 24) {real, imag} */,
  {32'hc2478511, 32'hc2300a7a} /* (7, 25, 23) {real, imag} */,
  {32'h402ddea8, 32'h4201d1d5} /* (7, 25, 22) {real, imag} */,
  {32'hc14e7c3a, 32'h420f2556} /* (7, 25, 21) {real, imag} */,
  {32'hc15acfde, 32'hc32254f5} /* (7, 25, 20) {real, imag} */,
  {32'h41e65905, 32'h42e66013} /* (7, 25, 19) {real, imag} */,
  {32'hc2dff83e, 32'hc2a5b1d5} /* (7, 25, 18) {real, imag} */,
  {32'hc1220340, 32'h4184ebc4} /* (7, 25, 17) {real, imag} */,
  {32'hc0d87890, 32'h00000000} /* (7, 25, 16) {real, imag} */,
  {32'hc1220340, 32'hc184ebc4} /* (7, 25, 15) {real, imag} */,
  {32'hc2dff83e, 32'h42a5b1d5} /* (7, 25, 14) {real, imag} */,
  {32'h41e65905, 32'hc2e66013} /* (7, 25, 13) {real, imag} */,
  {32'hc15acfde, 32'h432254f5} /* (7, 25, 12) {real, imag} */,
  {32'hc14e7c3a, 32'hc20f2556} /* (7, 25, 11) {real, imag} */,
  {32'h402ddea8, 32'hc201d1d5} /* (7, 25, 10) {real, imag} */,
  {32'hc2478511, 32'h42300a7a} /* (7, 25, 9) {real, imag} */,
  {32'hc187c573, 32'hc216c24f} /* (7, 25, 8) {real, imag} */,
  {32'h416a8085, 32'h430f02cc} /* (7, 25, 7) {real, imag} */,
  {32'h41b92754, 32'h41b49783} /* (7, 25, 6) {real, imag} */,
  {32'hc34a75f3, 32'hc2e9cf4c} /* (7, 25, 5) {real, imag} */,
  {32'h4341f538, 32'h417e0be8} /* (7, 25, 4) {real, imag} */,
  {32'hc1b37b88, 32'h42f19597} /* (7, 25, 3) {real, imag} */,
  {32'hc4aa006c, 32'hc3532284} /* (7, 25, 2) {real, imag} */,
  {32'h4552f8ef, 32'h440d4b01} /* (7, 25, 1) {real, imag} */,
  {32'h456cb6e8, 32'h00000000} /* (7, 25, 0) {real, imag} */,
  {32'h453e5a3c, 32'hc40cd597} /* (7, 24, 31) {real, imag} */,
  {32'hc4a5062a, 32'h43894126} /* (7, 24, 30) {real, imag} */,
  {32'hc0947940, 32'hc2ccac0b} /* (7, 24, 29) {real, imag} */,
  {32'h435304f9, 32'h41bcc8d4} /* (7, 24, 28) {real, imag} */,
  {32'hc376e830, 32'h42b75c64} /* (7, 24, 27) {real, imag} */,
  {32'hc23f0673, 32'hc1c92ea0} /* (7, 24, 26) {real, imag} */,
  {32'h41b95561, 32'hc2921ff0} /* (7, 24, 25) {real, imag} */,
  {32'hc2da6491, 32'hc205d5fc} /* (7, 24, 24) {real, imag} */,
  {32'hc0177ad0, 32'h410945a8} /* (7, 24, 23) {real, imag} */,
  {32'hc262c36c, 32'hc311474e} /* (7, 24, 22) {real, imag} */,
  {32'hc17cf000, 32'hc100bbde} /* (7, 24, 21) {real, imag} */,
  {32'hc15e6c6e, 32'h432c8900} /* (7, 24, 20) {real, imag} */,
  {32'hc22ac1bb, 32'hc2d8ae27} /* (7, 24, 19) {real, imag} */,
  {32'h42c16f9f, 32'h42305ab0} /* (7, 24, 18) {real, imag} */,
  {32'h40c5da5e, 32'hc1c03034} /* (7, 24, 17) {real, imag} */,
  {32'hc18ccc17, 32'h00000000} /* (7, 24, 16) {real, imag} */,
  {32'h40c5da5e, 32'h41c03034} /* (7, 24, 15) {real, imag} */,
  {32'h42c16f9f, 32'hc2305ab0} /* (7, 24, 14) {real, imag} */,
  {32'hc22ac1bb, 32'h42d8ae27} /* (7, 24, 13) {real, imag} */,
  {32'hc15e6c6e, 32'hc32c8900} /* (7, 24, 12) {real, imag} */,
  {32'hc17cf000, 32'h4100bbde} /* (7, 24, 11) {real, imag} */,
  {32'hc262c36c, 32'h4311474e} /* (7, 24, 10) {real, imag} */,
  {32'hc0177ad0, 32'hc10945a8} /* (7, 24, 9) {real, imag} */,
  {32'hc2da6491, 32'h4205d5fc} /* (7, 24, 8) {real, imag} */,
  {32'h41b95561, 32'h42921ff0} /* (7, 24, 7) {real, imag} */,
  {32'hc23f0673, 32'h41c92ea0} /* (7, 24, 6) {real, imag} */,
  {32'hc376e830, 32'hc2b75c64} /* (7, 24, 5) {real, imag} */,
  {32'h435304f9, 32'hc1bcc8d4} /* (7, 24, 4) {real, imag} */,
  {32'hc0947940, 32'h42ccac0b} /* (7, 24, 3) {real, imag} */,
  {32'hc4a5062a, 32'hc3894126} /* (7, 24, 2) {real, imag} */,
  {32'h453e5a3c, 32'h440cd597} /* (7, 24, 1) {real, imag} */,
  {32'h455728b6, 32'h00000000} /* (7, 24, 0) {real, imag} */,
  {32'h451615f4, 32'hc3dffe5a} /* (7, 23, 31) {real, imag} */,
  {32'hc48b8830, 32'h435403ee} /* (7, 23, 30) {real, imag} */,
  {32'hc337449a, 32'hc32a93d2} /* (7, 23, 29) {real, imag} */,
  {32'h42e3b5ba, 32'hc1ff1904} /* (7, 23, 28) {real, imag} */,
  {32'hc3025bdf, 32'h4297ef0a} /* (7, 23, 27) {real, imag} */,
  {32'h42cda87b, 32'h419c31a2} /* (7, 23, 26) {real, imag} */,
  {32'hc135771c, 32'hc0b64912} /* (7, 23, 25) {real, imag} */,
  {32'hc29e7f8d, 32'hc2119360} /* (7, 23, 24) {real, imag} */,
  {32'hc289866f, 32'h4288b392} /* (7, 23, 23) {real, imag} */,
  {32'hc1fa7dc2, 32'hc2024b2f} /* (7, 23, 22) {real, imag} */,
  {32'h4283a163, 32'h4156b792} /* (7, 23, 21) {real, imag} */,
  {32'h41a3aacd, 32'h4233dac8} /* (7, 23, 20) {real, imag} */,
  {32'h404562d8, 32'hc13813c2} /* (7, 23, 19) {real, imag} */,
  {32'h41ed6a9a, 32'h4191dd31} /* (7, 23, 18) {real, imag} */,
  {32'hc13fb4a2, 32'hc229c6e0} /* (7, 23, 17) {real, imag} */,
  {32'hc09abfdc, 32'h00000000} /* (7, 23, 16) {real, imag} */,
  {32'hc13fb4a2, 32'h4229c6e0} /* (7, 23, 15) {real, imag} */,
  {32'h41ed6a9a, 32'hc191dd31} /* (7, 23, 14) {real, imag} */,
  {32'h404562d8, 32'h413813c2} /* (7, 23, 13) {real, imag} */,
  {32'h41a3aacd, 32'hc233dac8} /* (7, 23, 12) {real, imag} */,
  {32'h4283a163, 32'hc156b792} /* (7, 23, 11) {real, imag} */,
  {32'hc1fa7dc2, 32'h42024b2f} /* (7, 23, 10) {real, imag} */,
  {32'hc289866f, 32'hc288b392} /* (7, 23, 9) {real, imag} */,
  {32'hc29e7f8d, 32'h42119360} /* (7, 23, 8) {real, imag} */,
  {32'hc135771c, 32'h40b64912} /* (7, 23, 7) {real, imag} */,
  {32'h42cda87b, 32'hc19c31a2} /* (7, 23, 6) {real, imag} */,
  {32'hc3025bdf, 32'hc297ef0a} /* (7, 23, 5) {real, imag} */,
  {32'h42e3b5ba, 32'h41ff1904} /* (7, 23, 4) {real, imag} */,
  {32'hc337449a, 32'h432a93d2} /* (7, 23, 3) {real, imag} */,
  {32'hc48b8830, 32'hc35403ee} /* (7, 23, 2) {real, imag} */,
  {32'h451615f4, 32'h43dffe5a} /* (7, 23, 1) {real, imag} */,
  {32'h4539a5ac, 32'h00000000} /* (7, 23, 0) {real, imag} */,
  {32'h44c5234c, 32'hc39ed4b8} /* (7, 22, 31) {real, imag} */,
  {32'hc46db420, 32'h431a86c0} /* (7, 22, 30) {real, imag} */,
  {32'hc34eb3a0, 32'hc35382fa} /* (7, 22, 29) {real, imag} */,
  {32'h430d5be6, 32'hc1de9d36} /* (7, 22, 28) {real, imag} */,
  {32'hc31bf16d, 32'h4324122b} /* (7, 22, 27) {real, imag} */,
  {32'h3fc6ab00, 32'h42955aca} /* (7, 22, 26) {real, imag} */,
  {32'h42afc747, 32'hc280da0a} /* (7, 22, 25) {real, imag} */,
  {32'hc2e22e2e, 32'h4057fa90} /* (7, 22, 24) {real, imag} */,
  {32'h424cfb04, 32'h3d404800} /* (7, 22, 23) {real, imag} */,
  {32'hc2ca76a7, 32'hc2473338} /* (7, 22, 22) {real, imag} */,
  {32'hc1d038e0, 32'hc26be4b2} /* (7, 22, 21) {real, imag} */,
  {32'h40a36798, 32'hc28904d5} /* (7, 22, 20) {real, imag} */,
  {32'h431c96e5, 32'h42844691} /* (7, 22, 19) {real, imag} */,
  {32'hc21e80e6, 32'hc29b7893} /* (7, 22, 18) {real, imag} */,
  {32'h3e54d780, 32'hc0c97988} /* (7, 22, 17) {real, imag} */,
  {32'hc0af4cda, 32'h00000000} /* (7, 22, 16) {real, imag} */,
  {32'h3e54d780, 32'h40c97988} /* (7, 22, 15) {real, imag} */,
  {32'hc21e80e6, 32'h429b7893} /* (7, 22, 14) {real, imag} */,
  {32'h431c96e5, 32'hc2844691} /* (7, 22, 13) {real, imag} */,
  {32'h40a36798, 32'h428904d5} /* (7, 22, 12) {real, imag} */,
  {32'hc1d038e0, 32'h426be4b2} /* (7, 22, 11) {real, imag} */,
  {32'hc2ca76a7, 32'h42473338} /* (7, 22, 10) {real, imag} */,
  {32'h424cfb04, 32'hbd404800} /* (7, 22, 9) {real, imag} */,
  {32'hc2e22e2e, 32'hc057fa90} /* (7, 22, 8) {real, imag} */,
  {32'h42afc747, 32'h4280da0a} /* (7, 22, 7) {real, imag} */,
  {32'h3fc6ab00, 32'hc2955aca} /* (7, 22, 6) {real, imag} */,
  {32'hc31bf16d, 32'hc324122b} /* (7, 22, 5) {real, imag} */,
  {32'h430d5be6, 32'h41de9d36} /* (7, 22, 4) {real, imag} */,
  {32'hc34eb3a0, 32'h435382fa} /* (7, 22, 3) {real, imag} */,
  {32'hc46db420, 32'hc31a86c0} /* (7, 22, 2) {real, imag} */,
  {32'h44c5234c, 32'h439ed4b8} /* (7, 22, 1) {real, imag} */,
  {32'h450d3684, 32'h00000000} /* (7, 22, 0) {real, imag} */,
  {32'h43e38668, 32'hc3442e3e} /* (7, 21, 31) {real, imag} */,
  {32'hc3993d1b, 32'hc33ea792} /* (7, 21, 30) {real, imag} */,
  {32'hc2eed2ed, 32'hc30d0030} /* (7, 21, 29) {real, imag} */,
  {32'h42df90a3, 32'h4279cd54} /* (7, 21, 28) {real, imag} */,
  {32'hc30414d0, 32'h42ff32e4} /* (7, 21, 27) {real, imag} */,
  {32'hc132da22, 32'h42605948} /* (7, 21, 26) {real, imag} */,
  {32'h423d21d0, 32'hc2d255fa} /* (7, 21, 25) {real, imag} */,
  {32'hc2923c1a, 32'hc2759ad7} /* (7, 21, 24) {real, imag} */,
  {32'hc224d22e, 32'h3ff0b328} /* (7, 21, 23) {real, imag} */,
  {32'h4211f378, 32'h425d0e27} /* (7, 21, 22) {real, imag} */,
  {32'hc2bcd9bc, 32'h426d7de1} /* (7, 21, 21) {real, imag} */,
  {32'h42260fb0, 32'h41b36750} /* (7, 21, 20) {real, imag} */,
  {32'hc17df13c, 32'h4203fab4} /* (7, 21, 19) {real, imag} */,
  {32'h42d41fae, 32'hc1e1427a} /* (7, 21, 18) {real, imag} */,
  {32'h4201ae96, 32'hc1f30e64} /* (7, 21, 17) {real, imag} */,
  {32'hc2bd2f0d, 32'h00000000} /* (7, 21, 16) {real, imag} */,
  {32'h4201ae96, 32'h41f30e64} /* (7, 21, 15) {real, imag} */,
  {32'h42d41fae, 32'h41e1427a} /* (7, 21, 14) {real, imag} */,
  {32'hc17df13c, 32'hc203fab4} /* (7, 21, 13) {real, imag} */,
  {32'h42260fb0, 32'hc1b36750} /* (7, 21, 12) {real, imag} */,
  {32'hc2bcd9bc, 32'hc26d7de1} /* (7, 21, 11) {real, imag} */,
  {32'h4211f378, 32'hc25d0e27} /* (7, 21, 10) {real, imag} */,
  {32'hc224d22e, 32'hbff0b328} /* (7, 21, 9) {real, imag} */,
  {32'hc2923c1a, 32'h42759ad7} /* (7, 21, 8) {real, imag} */,
  {32'h423d21d0, 32'h42d255fa} /* (7, 21, 7) {real, imag} */,
  {32'hc132da22, 32'hc2605948} /* (7, 21, 6) {real, imag} */,
  {32'hc30414d0, 32'hc2ff32e4} /* (7, 21, 5) {real, imag} */,
  {32'h42df90a3, 32'hc279cd54} /* (7, 21, 4) {real, imag} */,
  {32'hc2eed2ed, 32'h430d0030} /* (7, 21, 3) {real, imag} */,
  {32'hc3993d1b, 32'h433ea792} /* (7, 21, 2) {real, imag} */,
  {32'h43e38668, 32'h43442e3e} /* (7, 21, 1) {real, imag} */,
  {32'h449be120, 32'h00000000} /* (7, 21, 0) {real, imag} */,
  {32'hc4828468, 32'hc0f4bc80} /* (7, 20, 31) {real, imag} */,
  {32'h43f964bc, 32'hc3aad63d} /* (7, 20, 30) {real, imag} */,
  {32'hc31f2986, 32'hc2f38038} /* (7, 20, 29) {real, imag} */,
  {32'hc3006c99, 32'h42bd086b} /* (7, 20, 28) {real, imag} */,
  {32'h43399d10, 32'hc2bc72c8} /* (7, 20, 27) {real, imag} */,
  {32'h41dcd04e, 32'hc240d529} /* (7, 20, 26) {real, imag} */,
  {32'h421677a8, 32'hc19175b8} /* (7, 20, 25) {real, imag} */,
  {32'h40828ec8, 32'hc1c445cc} /* (7, 20, 24) {real, imag} */,
  {32'h420df310, 32'hc229b2b6} /* (7, 20, 23) {real, imag} */,
  {32'hc30e09d6, 32'h412f7444} /* (7, 20, 22) {real, imag} */,
  {32'hc250de3c, 32'hc1713562} /* (7, 20, 21) {real, imag} */,
  {32'hc1971ab4, 32'hc1b143c2} /* (7, 20, 20) {real, imag} */,
  {32'h40399690, 32'hc1e8863f} /* (7, 20, 19) {real, imag} */,
  {32'h42c3e7ce, 32'h42186284} /* (7, 20, 18) {real, imag} */,
  {32'h41458735, 32'hc1322812} /* (7, 20, 17) {real, imag} */,
  {32'h422f06c7, 32'h00000000} /* (7, 20, 16) {real, imag} */,
  {32'h41458735, 32'h41322812} /* (7, 20, 15) {real, imag} */,
  {32'h42c3e7ce, 32'hc2186284} /* (7, 20, 14) {real, imag} */,
  {32'h40399690, 32'h41e8863f} /* (7, 20, 13) {real, imag} */,
  {32'hc1971ab4, 32'h41b143c2} /* (7, 20, 12) {real, imag} */,
  {32'hc250de3c, 32'h41713562} /* (7, 20, 11) {real, imag} */,
  {32'hc30e09d6, 32'hc12f7444} /* (7, 20, 10) {real, imag} */,
  {32'h420df310, 32'h4229b2b6} /* (7, 20, 9) {real, imag} */,
  {32'h40828ec8, 32'h41c445cc} /* (7, 20, 8) {real, imag} */,
  {32'h421677a8, 32'h419175b8} /* (7, 20, 7) {real, imag} */,
  {32'h41dcd04e, 32'h4240d529} /* (7, 20, 6) {real, imag} */,
  {32'h43399d10, 32'h42bc72c8} /* (7, 20, 5) {real, imag} */,
  {32'hc3006c99, 32'hc2bd086b} /* (7, 20, 4) {real, imag} */,
  {32'hc31f2986, 32'h42f38038} /* (7, 20, 3) {real, imag} */,
  {32'h43f964bc, 32'h43aad63d} /* (7, 20, 2) {real, imag} */,
  {32'hc4828468, 32'h40f4bc80} /* (7, 20, 1) {real, imag} */,
  {32'hc39662c2, 32'h00000000} /* (7, 20, 0) {real, imag} */,
  {32'hc50413f1, 32'h430355e8} /* (7, 19, 31) {real, imag} */,
  {32'h447ae556, 32'hc3948bc9} /* (7, 19, 30) {real, imag} */,
  {32'hc378a950, 32'hc2ea6319} /* (7, 19, 29) {real, imag} */,
  {32'hc3233889, 32'hc261a246} /* (7, 19, 28) {real, imag} */,
  {32'h434910c9, 32'hc2ebb60c} /* (7, 19, 27) {real, imag} */,
  {32'h420ddc60, 32'hc163666d} /* (7, 19, 26) {real, imag} */,
  {32'hc22eba4d, 32'h4274ca4c} /* (7, 19, 25) {real, imag} */,
  {32'h400c0f68, 32'h419a073c} /* (7, 19, 24) {real, imag} */,
  {32'hc0224b90, 32'hc2c84baa} /* (7, 19, 23) {real, imag} */,
  {32'hc1f2b706, 32'hc1b1a0a6} /* (7, 19, 22) {real, imag} */,
  {32'h42b155e5, 32'h4286252c} /* (7, 19, 21) {real, imag} */,
  {32'h416abc52, 32'h421f471e} /* (7, 19, 20) {real, imag} */,
  {32'hc18617d0, 32'hc295c002} /* (7, 19, 19) {real, imag} */,
  {32'h42a1b958, 32'hc2169c82} /* (7, 19, 18) {real, imag} */,
  {32'h40ad6bcd, 32'h425e07e8} /* (7, 19, 17) {real, imag} */,
  {32'hc2cebd75, 32'h00000000} /* (7, 19, 16) {real, imag} */,
  {32'h40ad6bcd, 32'hc25e07e8} /* (7, 19, 15) {real, imag} */,
  {32'h42a1b958, 32'h42169c82} /* (7, 19, 14) {real, imag} */,
  {32'hc18617d0, 32'h4295c002} /* (7, 19, 13) {real, imag} */,
  {32'h416abc52, 32'hc21f471e} /* (7, 19, 12) {real, imag} */,
  {32'h42b155e5, 32'hc286252c} /* (7, 19, 11) {real, imag} */,
  {32'hc1f2b706, 32'h41b1a0a6} /* (7, 19, 10) {real, imag} */,
  {32'hc0224b90, 32'h42c84baa} /* (7, 19, 9) {real, imag} */,
  {32'h400c0f68, 32'hc19a073c} /* (7, 19, 8) {real, imag} */,
  {32'hc22eba4d, 32'hc274ca4c} /* (7, 19, 7) {real, imag} */,
  {32'h420ddc60, 32'h4163666d} /* (7, 19, 6) {real, imag} */,
  {32'h434910c9, 32'h42ebb60c} /* (7, 19, 5) {real, imag} */,
  {32'hc3233889, 32'h4261a246} /* (7, 19, 4) {real, imag} */,
  {32'hc378a950, 32'h42ea6319} /* (7, 19, 3) {real, imag} */,
  {32'h447ae556, 32'h43948bc9} /* (7, 19, 2) {real, imag} */,
  {32'hc50413f1, 32'hc30355e8} /* (7, 19, 1) {real, imag} */,
  {32'hc47730ad, 32'h00000000} /* (7, 19, 0) {real, imag} */,
  {32'hc5332d74, 32'h4387144d} /* (7, 18, 31) {real, imag} */,
  {32'h44925f32, 32'hc39a345a} /* (7, 18, 30) {real, imag} */,
  {32'hc339f1dc, 32'hc202e0cd} /* (7, 18, 29) {real, imag} */,
  {32'hc2e6ab1b, 32'hc18dc118} /* (7, 18, 28) {real, imag} */,
  {32'h42d87f34, 32'hc0d3c380} /* (7, 18, 27) {real, imag} */,
  {32'h4315d629, 32'h416c8256} /* (7, 18, 26) {real, imag} */,
  {32'hc283cbac, 32'h40780dac} /* (7, 18, 25) {real, imag} */,
  {32'h4219a0be, 32'h424c5edf} /* (7, 18, 24) {real, imag} */,
  {32'h42681c90, 32'hc2edcfbe} /* (7, 18, 23) {real, imag} */,
  {32'h4216de82, 32'h42d590dc} /* (7, 18, 22) {real, imag} */,
  {32'hc2254cb8, 32'hc342ec8f} /* (7, 18, 21) {real, imag} */,
  {32'hc2003f76, 32'h4101dbac} /* (7, 18, 20) {real, imag} */,
  {32'hc1402f5a, 32'hc2647d76} /* (7, 18, 19) {real, imag} */,
  {32'h40e5f51c, 32'hc0c1b570} /* (7, 18, 18) {real, imag} */,
  {32'h41919d0e, 32'hc13975d4} /* (7, 18, 17) {real, imag} */,
  {32'hc23e2680, 32'h00000000} /* (7, 18, 16) {real, imag} */,
  {32'h41919d0e, 32'h413975d4} /* (7, 18, 15) {real, imag} */,
  {32'h40e5f51c, 32'h40c1b570} /* (7, 18, 14) {real, imag} */,
  {32'hc1402f5a, 32'h42647d76} /* (7, 18, 13) {real, imag} */,
  {32'hc2003f76, 32'hc101dbac} /* (7, 18, 12) {real, imag} */,
  {32'hc2254cb8, 32'h4342ec8f} /* (7, 18, 11) {real, imag} */,
  {32'h4216de82, 32'hc2d590dc} /* (7, 18, 10) {real, imag} */,
  {32'h42681c90, 32'h42edcfbe} /* (7, 18, 9) {real, imag} */,
  {32'h4219a0be, 32'hc24c5edf} /* (7, 18, 8) {real, imag} */,
  {32'hc283cbac, 32'hc0780dac} /* (7, 18, 7) {real, imag} */,
  {32'h4315d629, 32'hc16c8256} /* (7, 18, 6) {real, imag} */,
  {32'h42d87f34, 32'h40d3c380} /* (7, 18, 5) {real, imag} */,
  {32'hc2e6ab1b, 32'h418dc118} /* (7, 18, 4) {real, imag} */,
  {32'hc339f1dc, 32'h4202e0cd} /* (7, 18, 3) {real, imag} */,
  {32'h44925f32, 32'h439a345a} /* (7, 18, 2) {real, imag} */,
  {32'hc5332d74, 32'hc387144d} /* (7, 18, 1) {real, imag} */,
  {32'hc4cd2b7f, 32'h00000000} /* (7, 18, 0) {real, imag} */,
  {32'hc549cf34, 32'h4393a56d} /* (7, 17, 31) {real, imag} */,
  {32'h44919d4a, 32'hc39f6a7e} /* (7, 17, 30) {real, imag} */,
  {32'hc2741a9c, 32'hc2372b08} /* (7, 17, 29) {real, imag} */,
  {32'hc324bf63, 32'hc1ebeb36} /* (7, 17, 28) {real, imag} */,
  {32'h435837d6, 32'h42a348ae} /* (7, 17, 27) {real, imag} */,
  {32'h42b5cc6c, 32'h426c9fe5} /* (7, 17, 26) {real, imag} */,
  {32'h429b8e89, 32'h4238e983} /* (7, 17, 25) {real, imag} */,
  {32'h4224891b, 32'hc2242e3f} /* (7, 17, 24) {real, imag} */,
  {32'h429d6d7d, 32'h430276aa} /* (7, 17, 23) {real, imag} */,
  {32'h413f56d6, 32'hc1ec7159} /* (7, 17, 22) {real, imag} */,
  {32'h42948902, 32'hc2c6ea42} /* (7, 17, 21) {real, imag} */,
  {32'hc304631c, 32'hc230c80a} /* (7, 17, 20) {real, imag} */,
  {32'h40b08e42, 32'hc248f26c} /* (7, 17, 19) {real, imag} */,
  {32'hc018b218, 32'h42164830} /* (7, 17, 18) {real, imag} */,
  {32'h42026ed4, 32'hc0134cf0} /* (7, 17, 17) {real, imag} */,
  {32'hc1db1b78, 32'h00000000} /* (7, 17, 16) {real, imag} */,
  {32'h42026ed4, 32'h40134cf0} /* (7, 17, 15) {real, imag} */,
  {32'hc018b218, 32'hc2164830} /* (7, 17, 14) {real, imag} */,
  {32'h40b08e42, 32'h4248f26c} /* (7, 17, 13) {real, imag} */,
  {32'hc304631c, 32'h4230c80a} /* (7, 17, 12) {real, imag} */,
  {32'h42948902, 32'h42c6ea42} /* (7, 17, 11) {real, imag} */,
  {32'h413f56d6, 32'h41ec7159} /* (7, 17, 10) {real, imag} */,
  {32'h429d6d7d, 32'hc30276aa} /* (7, 17, 9) {real, imag} */,
  {32'h4224891b, 32'h42242e3f} /* (7, 17, 8) {real, imag} */,
  {32'h429b8e89, 32'hc238e983} /* (7, 17, 7) {real, imag} */,
  {32'h42b5cc6c, 32'hc26c9fe5} /* (7, 17, 6) {real, imag} */,
  {32'h435837d6, 32'hc2a348ae} /* (7, 17, 5) {real, imag} */,
  {32'hc324bf63, 32'h41ebeb36} /* (7, 17, 4) {real, imag} */,
  {32'hc2741a9c, 32'h42372b08} /* (7, 17, 3) {real, imag} */,
  {32'h44919d4a, 32'h439f6a7e} /* (7, 17, 2) {real, imag} */,
  {32'hc549cf34, 32'hc393a56d} /* (7, 17, 1) {real, imag} */,
  {32'hc50c5fad, 32'h00000000} /* (7, 17, 0) {real, imag} */,
  {32'hc5505974, 32'h4390c12e} /* (7, 16, 31) {real, imag} */,
  {32'h4498c566, 32'hc3158007} /* (7, 16, 30) {real, imag} */,
  {32'hc293f79b, 32'hc313a01b} /* (7, 16, 29) {real, imag} */,
  {32'hc3233d27, 32'h4283031d} /* (7, 16, 28) {real, imag} */,
  {32'h42ec9800, 32'hc2355008} /* (7, 16, 27) {real, imag} */,
  {32'h42364e96, 32'hc2ac5477} /* (7, 16, 26) {real, imag} */,
  {32'h42d18db2, 32'hc2a4fd44} /* (7, 16, 25) {real, imag} */,
  {32'h4295bb40, 32'hc29546eb} /* (7, 16, 24) {real, imag} */,
  {32'h42773028, 32'h42066969} /* (7, 16, 23) {real, imag} */,
  {32'hc1c9f1c3, 32'h428bbe1c} /* (7, 16, 22) {real, imag} */,
  {32'h42c67c44, 32'hc22adb1e} /* (7, 16, 21) {real, imag} */,
  {32'h4209e67f, 32'hc2b615be} /* (7, 16, 20) {real, imag} */,
  {32'hc2b4953a, 32'hc207478d} /* (7, 16, 19) {real, imag} */,
  {32'h410c26a8, 32'h41b328ee} /* (7, 16, 18) {real, imag} */,
  {32'hc13a7fb7, 32'h419c1dc5} /* (7, 16, 17) {real, imag} */,
  {32'hc2a7055e, 32'h00000000} /* (7, 16, 16) {real, imag} */,
  {32'hc13a7fb7, 32'hc19c1dc5} /* (7, 16, 15) {real, imag} */,
  {32'h410c26a8, 32'hc1b328ee} /* (7, 16, 14) {real, imag} */,
  {32'hc2b4953a, 32'h4207478d} /* (7, 16, 13) {real, imag} */,
  {32'h4209e67f, 32'h42b615be} /* (7, 16, 12) {real, imag} */,
  {32'h42c67c44, 32'h422adb1e} /* (7, 16, 11) {real, imag} */,
  {32'hc1c9f1c3, 32'hc28bbe1c} /* (7, 16, 10) {real, imag} */,
  {32'h42773028, 32'hc2066969} /* (7, 16, 9) {real, imag} */,
  {32'h4295bb40, 32'h429546eb} /* (7, 16, 8) {real, imag} */,
  {32'h42d18db2, 32'h42a4fd44} /* (7, 16, 7) {real, imag} */,
  {32'h42364e96, 32'h42ac5477} /* (7, 16, 6) {real, imag} */,
  {32'h42ec9800, 32'h42355008} /* (7, 16, 5) {real, imag} */,
  {32'hc3233d27, 32'hc283031d} /* (7, 16, 4) {real, imag} */,
  {32'hc293f79b, 32'h4313a01b} /* (7, 16, 3) {real, imag} */,
  {32'h4498c566, 32'h43158007} /* (7, 16, 2) {real, imag} */,
  {32'hc5505974, 32'hc390c12e} /* (7, 16, 1) {real, imag} */,
  {32'hc5197b68, 32'h00000000} /* (7, 16, 0) {real, imag} */,
  {32'hc553f368, 32'h43a9c467} /* (7, 15, 31) {real, imag} */,
  {32'h449e8c36, 32'hc2de9443} /* (7, 15, 30) {real, imag} */,
  {32'hc1176d30, 32'hc2d463cc} /* (7, 15, 29) {real, imag} */,
  {32'hc31bd419, 32'hc304a3af} /* (7, 15, 28) {real, imag} */,
  {32'h42f68160, 32'hc335d0d1} /* (7, 15, 27) {real, imag} */,
  {32'h42190144, 32'hc2d8b540} /* (7, 15, 26) {real, imag} */,
  {32'hc2a49f63, 32'hc265f4dd} /* (7, 15, 25) {real, imag} */,
  {32'h42f9e6cc, 32'hc2293335} /* (7, 15, 24) {real, imag} */,
  {32'hc2315bc6, 32'hc2fb2225} /* (7, 15, 23) {real, imag} */,
  {32'hc15e5a56, 32'h4226ec78} /* (7, 15, 22) {real, imag} */,
  {32'h41fcae10, 32'hc0976c28} /* (7, 15, 21) {real, imag} */,
  {32'h428b6378, 32'hc2bdc789} /* (7, 15, 20) {real, imag} */,
  {32'h4209bd06, 32'h42373384} /* (7, 15, 19) {real, imag} */,
  {32'h42119c24, 32'h424097fc} /* (7, 15, 18) {real, imag} */,
  {32'h42238870, 32'hc25bbe63} /* (7, 15, 17) {real, imag} */,
  {32'h413e0b90, 32'h00000000} /* (7, 15, 16) {real, imag} */,
  {32'h42238870, 32'h425bbe63} /* (7, 15, 15) {real, imag} */,
  {32'h42119c24, 32'hc24097fc} /* (7, 15, 14) {real, imag} */,
  {32'h4209bd06, 32'hc2373384} /* (7, 15, 13) {real, imag} */,
  {32'h428b6378, 32'h42bdc789} /* (7, 15, 12) {real, imag} */,
  {32'h41fcae10, 32'h40976c28} /* (7, 15, 11) {real, imag} */,
  {32'hc15e5a56, 32'hc226ec78} /* (7, 15, 10) {real, imag} */,
  {32'hc2315bc6, 32'h42fb2225} /* (7, 15, 9) {real, imag} */,
  {32'h42f9e6cc, 32'h42293335} /* (7, 15, 8) {real, imag} */,
  {32'hc2a49f63, 32'h4265f4dd} /* (7, 15, 7) {real, imag} */,
  {32'h42190144, 32'h42d8b540} /* (7, 15, 6) {real, imag} */,
  {32'h42f68160, 32'h4335d0d1} /* (7, 15, 5) {real, imag} */,
  {32'hc31bd419, 32'h4304a3af} /* (7, 15, 4) {real, imag} */,
  {32'hc1176d30, 32'h42d463cc} /* (7, 15, 3) {real, imag} */,
  {32'h449e8c36, 32'h42de9443} /* (7, 15, 2) {real, imag} */,
  {32'hc553f368, 32'hc3a9c467} /* (7, 15, 1) {real, imag} */,
  {32'hc5265e19, 32'h00000000} /* (7, 15, 0) {real, imag} */,
  {32'hc53b27fc, 32'h42fd296c} /* (7, 14, 31) {real, imag} */,
  {32'h449d6130, 32'hc3763dd0} /* (7, 14, 30) {real, imag} */,
  {32'h426ebc26, 32'h4184287a} /* (7, 14, 29) {real, imag} */,
  {32'hc34c12ba, 32'hc2e061d0} /* (7, 14, 28) {real, imag} */,
  {32'h4302ba9b, 32'hc2d03ede} /* (7, 14, 27) {real, imag} */,
  {32'h4286d5d2, 32'hc25dee3e} /* (7, 14, 26) {real, imag} */,
  {32'hc235ee4c, 32'h41d58690} /* (7, 14, 25) {real, imag} */,
  {32'h4103c7c6, 32'hc1c3cee2} /* (7, 14, 24) {real, imag} */,
  {32'hc2ae5360, 32'hc1647700} /* (7, 14, 23) {real, imag} */,
  {32'h42888a1b, 32'hc232c840} /* (7, 14, 22) {real, imag} */,
  {32'h42962e15, 32'hc19e2db8} /* (7, 14, 21) {real, imag} */,
  {32'h42608ac2, 32'hc2abfbe2} /* (7, 14, 20) {real, imag} */,
  {32'h421df9a6, 32'h40f87be0} /* (7, 14, 19) {real, imag} */,
  {32'hc2660df0, 32'hc240a1f4} /* (7, 14, 18) {real, imag} */,
  {32'h426c4569, 32'h421c87fe} /* (7, 14, 17) {real, imag} */,
  {32'h42de0812, 32'h00000000} /* (7, 14, 16) {real, imag} */,
  {32'h426c4569, 32'hc21c87fe} /* (7, 14, 15) {real, imag} */,
  {32'hc2660df0, 32'h4240a1f4} /* (7, 14, 14) {real, imag} */,
  {32'h421df9a6, 32'hc0f87be0} /* (7, 14, 13) {real, imag} */,
  {32'h42608ac2, 32'h42abfbe2} /* (7, 14, 12) {real, imag} */,
  {32'h42962e15, 32'h419e2db8} /* (7, 14, 11) {real, imag} */,
  {32'h42888a1b, 32'h4232c840} /* (7, 14, 10) {real, imag} */,
  {32'hc2ae5360, 32'h41647700} /* (7, 14, 9) {real, imag} */,
  {32'h4103c7c6, 32'h41c3cee2} /* (7, 14, 8) {real, imag} */,
  {32'hc235ee4c, 32'hc1d58690} /* (7, 14, 7) {real, imag} */,
  {32'h4286d5d2, 32'h425dee3e} /* (7, 14, 6) {real, imag} */,
  {32'h4302ba9b, 32'h42d03ede} /* (7, 14, 5) {real, imag} */,
  {32'hc34c12ba, 32'h42e061d0} /* (7, 14, 4) {real, imag} */,
  {32'h426ebc26, 32'hc184287a} /* (7, 14, 3) {real, imag} */,
  {32'h449d6130, 32'h43763dd0} /* (7, 14, 2) {real, imag} */,
  {32'hc53b27fc, 32'hc2fd296c} /* (7, 14, 1) {real, imag} */,
  {32'hc51f5728, 32'h00000000} /* (7, 14, 0) {real, imag} */,
  {32'hc51e1ab5, 32'h4109a200} /* (7, 13, 31) {real, imag} */,
  {32'h448c36a5, 32'hc310f7f6} /* (7, 13, 30) {real, imag} */,
  {32'h42227c7e, 32'hc24c774a} /* (7, 13, 29) {real, imag} */,
  {32'hc306e433, 32'h401615e0} /* (7, 13, 28) {real, imag} */,
  {32'h4361dd67, 32'hc2748a98} /* (7, 13, 27) {real, imag} */,
  {32'h4293c8bc, 32'h418975be} /* (7, 13, 26) {real, imag} */,
  {32'hc3130b55, 32'h42abe742} /* (7, 13, 25) {real, imag} */,
  {32'h4203474e, 32'hc320956a} /* (7, 13, 24) {real, imag} */,
  {32'h42e55b92, 32'hc18e4b4e} /* (7, 13, 23) {real, imag} */,
  {32'hc0db7a48, 32'h424774cf} /* (7, 13, 22) {real, imag} */,
  {32'hc27c53ca, 32'h418dda16} /* (7, 13, 21) {real, imag} */,
  {32'h41b6eceb, 32'hc270d65a} /* (7, 13, 20) {real, imag} */,
  {32'hc1920586, 32'hc12c9b18} /* (7, 13, 19) {real, imag} */,
  {32'h4183a464, 32'h4144d2f0} /* (7, 13, 18) {real, imag} */,
  {32'h410be1fe, 32'hc298aa40} /* (7, 13, 17) {real, imag} */,
  {32'h42a3c4ab, 32'h00000000} /* (7, 13, 16) {real, imag} */,
  {32'h410be1fe, 32'h4298aa40} /* (7, 13, 15) {real, imag} */,
  {32'h4183a464, 32'hc144d2f0} /* (7, 13, 14) {real, imag} */,
  {32'hc1920586, 32'h412c9b18} /* (7, 13, 13) {real, imag} */,
  {32'h41b6eceb, 32'h4270d65a} /* (7, 13, 12) {real, imag} */,
  {32'hc27c53ca, 32'hc18dda16} /* (7, 13, 11) {real, imag} */,
  {32'hc0db7a48, 32'hc24774cf} /* (7, 13, 10) {real, imag} */,
  {32'h42e55b92, 32'h418e4b4e} /* (7, 13, 9) {real, imag} */,
  {32'h4203474e, 32'h4320956a} /* (7, 13, 8) {real, imag} */,
  {32'hc3130b55, 32'hc2abe742} /* (7, 13, 7) {real, imag} */,
  {32'h4293c8bc, 32'hc18975be} /* (7, 13, 6) {real, imag} */,
  {32'h4361dd67, 32'h42748a98} /* (7, 13, 5) {real, imag} */,
  {32'hc306e433, 32'hc01615e0} /* (7, 13, 4) {real, imag} */,
  {32'h42227c7e, 32'h424c774a} /* (7, 13, 3) {real, imag} */,
  {32'h448c36a5, 32'h4310f7f6} /* (7, 13, 2) {real, imag} */,
  {32'hc51e1ab5, 32'hc109a200} /* (7, 13, 1) {real, imag} */,
  {32'hc5073d23, 32'h00000000} /* (7, 13, 0) {real, imag} */,
  {32'hc4e195a4, 32'h416daf40} /* (7, 12, 31) {real, imag} */,
  {32'h446f9e1c, 32'hc24fc0f8} /* (7, 12, 30) {real, imag} */,
  {32'h43951847, 32'h429c81e4} /* (7, 12, 29) {real, imag} */,
  {32'hc30e20a3, 32'hc248967a} /* (7, 12, 28) {real, imag} */,
  {32'h420db572, 32'hc14a7640} /* (7, 12, 27) {real, imag} */,
  {32'h42446cd1, 32'hc239ff35} /* (7, 12, 26) {real, imag} */,
  {32'hc2c2a158, 32'hc3224fcf} /* (7, 12, 25) {real, imag} */,
  {32'hc174d86c, 32'hc30b8d42} /* (7, 12, 24) {real, imag} */,
  {32'h3f1892a0, 32'h42731caa} /* (7, 12, 23) {real, imag} */,
  {32'hc207b78f, 32'h42a591ce} /* (7, 12, 22) {real, imag} */,
  {32'h422d8ae0, 32'hc244d710} /* (7, 12, 21) {real, imag} */,
  {32'h40f44a52, 32'hc29063a6} /* (7, 12, 20) {real, imag} */,
  {32'h428ba7b4, 32'h4206774a} /* (7, 12, 19) {real, imag} */,
  {32'hc22d2ff3, 32'hbfcbe4f0} /* (7, 12, 18) {real, imag} */,
  {32'hc179fee5, 32'h41c86843} /* (7, 12, 17) {real, imag} */,
  {32'hc198301e, 32'h00000000} /* (7, 12, 16) {real, imag} */,
  {32'hc179fee5, 32'hc1c86843} /* (7, 12, 15) {real, imag} */,
  {32'hc22d2ff3, 32'h3fcbe4f0} /* (7, 12, 14) {real, imag} */,
  {32'h428ba7b4, 32'hc206774a} /* (7, 12, 13) {real, imag} */,
  {32'h40f44a52, 32'h429063a6} /* (7, 12, 12) {real, imag} */,
  {32'h422d8ae0, 32'h4244d710} /* (7, 12, 11) {real, imag} */,
  {32'hc207b78f, 32'hc2a591ce} /* (7, 12, 10) {real, imag} */,
  {32'h3f1892a0, 32'hc2731caa} /* (7, 12, 9) {real, imag} */,
  {32'hc174d86c, 32'h430b8d42} /* (7, 12, 8) {real, imag} */,
  {32'hc2c2a158, 32'h43224fcf} /* (7, 12, 7) {real, imag} */,
  {32'h42446cd1, 32'h4239ff35} /* (7, 12, 6) {real, imag} */,
  {32'h420db572, 32'h414a7640} /* (7, 12, 5) {real, imag} */,
  {32'hc30e20a3, 32'h4248967a} /* (7, 12, 4) {real, imag} */,
  {32'h43951847, 32'hc29c81e4} /* (7, 12, 3) {real, imag} */,
  {32'h446f9e1c, 32'h424fc0f8} /* (7, 12, 2) {real, imag} */,
  {32'hc4e195a4, 32'hc16daf40} /* (7, 12, 1) {real, imag} */,
  {32'hc4be5c64, 32'h00000000} /* (7, 12, 0) {real, imag} */,
  {32'hc464e748, 32'hc380fdb5} /* (7, 11, 31) {real, imag} */,
  {32'h4400e71c, 32'hc2901873} /* (7, 11, 30) {real, imag} */,
  {32'h4330d081, 32'h42a989a3} /* (7, 11, 29) {real, imag} */,
  {32'hc32789b0, 32'hc2e08dce} /* (7, 11, 28) {real, imag} */,
  {32'h41813b60, 32'hc20f3d49} /* (7, 11, 27) {real, imag} */,
  {32'hc28e3941, 32'h41a694ef} /* (7, 11, 26) {real, imag} */,
  {32'hc25f1294, 32'hc247f0f0} /* (7, 11, 25) {real, imag} */,
  {32'h4303a5c3, 32'hc32326f7} /* (7, 11, 24) {real, imag} */,
  {32'hc1938fbf, 32'h41a78a4c} /* (7, 11, 23) {real, imag} */,
  {32'hc1c068a3, 32'h40f8a818} /* (7, 11, 22) {real, imag} */,
  {32'h42561bf5, 32'hc238f143} /* (7, 11, 21) {real, imag} */,
  {32'hc21e10a8, 32'hc20a8a5c} /* (7, 11, 20) {real, imag} */,
  {32'hc2d892be, 32'hc28ddf68} /* (7, 11, 19) {real, imag} */,
  {32'h4146ead0, 32'hc254f02f} /* (7, 11, 18) {real, imag} */,
  {32'h4060d150, 32'h42427b80} /* (7, 11, 17) {real, imag} */,
  {32'h4271f0e6, 32'h00000000} /* (7, 11, 16) {real, imag} */,
  {32'h4060d150, 32'hc2427b80} /* (7, 11, 15) {real, imag} */,
  {32'h4146ead0, 32'h4254f02f} /* (7, 11, 14) {real, imag} */,
  {32'hc2d892be, 32'h428ddf68} /* (7, 11, 13) {real, imag} */,
  {32'hc21e10a8, 32'h420a8a5c} /* (7, 11, 12) {real, imag} */,
  {32'h42561bf5, 32'h4238f143} /* (7, 11, 11) {real, imag} */,
  {32'hc1c068a3, 32'hc0f8a818} /* (7, 11, 10) {real, imag} */,
  {32'hc1938fbf, 32'hc1a78a4c} /* (7, 11, 9) {real, imag} */,
  {32'h4303a5c3, 32'h432326f7} /* (7, 11, 8) {real, imag} */,
  {32'hc25f1294, 32'h4247f0f0} /* (7, 11, 7) {real, imag} */,
  {32'hc28e3941, 32'hc1a694ef} /* (7, 11, 6) {real, imag} */,
  {32'h41813b60, 32'h420f3d49} /* (7, 11, 5) {real, imag} */,
  {32'hc32789b0, 32'h42e08dce} /* (7, 11, 4) {real, imag} */,
  {32'h4330d081, 32'hc2a989a3} /* (7, 11, 3) {real, imag} */,
  {32'h4400e71c, 32'h42901873} /* (7, 11, 2) {real, imag} */,
  {32'hc464e748, 32'h4380fdb5} /* (7, 11, 1) {real, imag} */,
  {32'hc3f6881e, 32'h00000000} /* (7, 11, 0) {real, imag} */,
  {32'h441e5e48, 32'hc410f856} /* (7, 10, 31) {real, imag} */,
  {32'hc378054a, 32'h4342b4d4} /* (7, 10, 30) {real, imag} */,
  {32'h430e95a4, 32'hc1a2d124} /* (7, 10, 29) {real, imag} */,
  {32'h4097e1d0, 32'hc30224a4} /* (7, 10, 28) {real, imag} */,
  {32'h42858e82, 32'h4294be94} /* (7, 10, 27) {real, imag} */,
  {32'hc2b29482, 32'h4183c408} /* (7, 10, 26) {real, imag} */,
  {32'h430ffbcc, 32'h41a16df9} /* (7, 10, 25) {real, imag} */,
  {32'hc24bffeb, 32'h418a43da} /* (7, 10, 24) {real, imag} */,
  {32'h41bcb0b0, 32'hc2df3d0a} /* (7, 10, 23) {real, imag} */,
  {32'hc220efee, 32'h40ce0da4} /* (7, 10, 22) {real, imag} */,
  {32'h3fb67a88, 32'h425df7f4} /* (7, 10, 21) {real, imag} */,
  {32'hc216beb5, 32'hc2bd9a1b} /* (7, 10, 20) {real, imag} */,
  {32'h42ab8612, 32'h41458d6a} /* (7, 10, 19) {real, imag} */,
  {32'hc0979a20, 32'h42256a30} /* (7, 10, 18) {real, imag} */,
  {32'h42008d66, 32'hc0b50f48} /* (7, 10, 17) {real, imag} */,
  {32'hc198bb92, 32'h00000000} /* (7, 10, 16) {real, imag} */,
  {32'h42008d66, 32'h40b50f48} /* (7, 10, 15) {real, imag} */,
  {32'hc0979a20, 32'hc2256a30} /* (7, 10, 14) {real, imag} */,
  {32'h42ab8612, 32'hc1458d6a} /* (7, 10, 13) {real, imag} */,
  {32'hc216beb5, 32'h42bd9a1b} /* (7, 10, 12) {real, imag} */,
  {32'h3fb67a88, 32'hc25df7f4} /* (7, 10, 11) {real, imag} */,
  {32'hc220efee, 32'hc0ce0da4} /* (7, 10, 10) {real, imag} */,
  {32'h41bcb0b0, 32'h42df3d0a} /* (7, 10, 9) {real, imag} */,
  {32'hc24bffeb, 32'hc18a43da} /* (7, 10, 8) {real, imag} */,
  {32'h430ffbcc, 32'hc1a16df9} /* (7, 10, 7) {real, imag} */,
  {32'hc2b29482, 32'hc183c408} /* (7, 10, 6) {real, imag} */,
  {32'h42858e82, 32'hc294be94} /* (7, 10, 5) {real, imag} */,
  {32'h4097e1d0, 32'h430224a4} /* (7, 10, 4) {real, imag} */,
  {32'h430e95a4, 32'h41a2d124} /* (7, 10, 3) {real, imag} */,
  {32'hc378054a, 32'hc342b4d4} /* (7, 10, 2) {real, imag} */,
  {32'h441e5e48, 32'h4410f856} /* (7, 10, 1) {real, imag} */,
  {32'h442e2e40, 32'h00000000} /* (7, 10, 0) {real, imag} */,
  {32'h44d51beb, 32'hc469e8dd} /* (7, 9, 31) {real, imag} */,
  {32'hc427d1aa, 32'h43c91f53} /* (7, 9, 30) {real, imag} */,
  {32'h438fc30e, 32'h42a17e23} /* (7, 9, 29) {real, imag} */,
  {32'h431cb173, 32'hc34c04be} /* (7, 9, 28) {real, imag} */,
  {32'h3f7ea100, 32'h4336f827} /* (7, 9, 27) {real, imag} */,
  {32'hc29d4a23, 32'hc0cbaff2} /* (7, 9, 26) {real, imag} */,
  {32'hc26bde71, 32'h418af294} /* (7, 9, 25) {real, imag} */,
  {32'hc24432c6, 32'hc0f91134} /* (7, 9, 24) {real, imag} */,
  {32'h42ea5aa5, 32'h41055b18} /* (7, 9, 23) {real, imag} */,
  {32'hc2d4a7de, 32'hc1f41596} /* (7, 9, 22) {real, imag} */,
  {32'hc2a705d5, 32'h41df1dcf} /* (7, 9, 21) {real, imag} */,
  {32'h408bc9d4, 32'h4293b578} /* (7, 9, 20) {real, imag} */,
  {32'h416e64da, 32'hc119b566} /* (7, 9, 19) {real, imag} */,
  {32'hc18e301e, 32'h4299fc66} /* (7, 9, 18) {real, imag} */,
  {32'hc25bbe38, 32'hc19d48b3} /* (7, 9, 17) {real, imag} */,
  {32'hc127b3b8, 32'h00000000} /* (7, 9, 16) {real, imag} */,
  {32'hc25bbe38, 32'h419d48b3} /* (7, 9, 15) {real, imag} */,
  {32'hc18e301e, 32'hc299fc66} /* (7, 9, 14) {real, imag} */,
  {32'h416e64da, 32'h4119b566} /* (7, 9, 13) {real, imag} */,
  {32'h408bc9d4, 32'hc293b578} /* (7, 9, 12) {real, imag} */,
  {32'hc2a705d5, 32'hc1df1dcf} /* (7, 9, 11) {real, imag} */,
  {32'hc2d4a7de, 32'h41f41596} /* (7, 9, 10) {real, imag} */,
  {32'h42ea5aa5, 32'hc1055b18} /* (7, 9, 9) {real, imag} */,
  {32'hc24432c6, 32'h40f91134} /* (7, 9, 8) {real, imag} */,
  {32'hc26bde71, 32'hc18af294} /* (7, 9, 7) {real, imag} */,
  {32'hc29d4a23, 32'h40cbaff2} /* (7, 9, 6) {real, imag} */,
  {32'h3f7ea100, 32'hc336f827} /* (7, 9, 5) {real, imag} */,
  {32'h431cb173, 32'h434c04be} /* (7, 9, 4) {real, imag} */,
  {32'h438fc30e, 32'hc2a17e23} /* (7, 9, 3) {real, imag} */,
  {32'hc427d1aa, 32'hc3c91f53} /* (7, 9, 2) {real, imag} */,
  {32'h44d51beb, 32'h4469e8dd} /* (7, 9, 1) {real, imag} */,
  {32'h44fd1d40, 32'h00000000} /* (7, 9, 0) {real, imag} */,
  {32'h450f6040, 32'hc485f3d4} /* (7, 8, 31) {real, imag} */,
  {32'hc443b66b, 32'h43e2279e} /* (7, 8, 30) {real, imag} */,
  {32'h434067a8, 32'h430ff5c6} /* (7, 8, 29) {real, imag} */,
  {32'h4330a681, 32'hc321128a} /* (7, 8, 28) {real, imag} */,
  {32'hc33613fa, 32'h43114998} /* (7, 8, 27) {real, imag} */,
  {32'hc1aa397e, 32'h429df706} /* (7, 8, 26) {real, imag} */,
  {32'h416702fa, 32'hc229cdbc} /* (7, 8, 25) {real, imag} */,
  {32'hc1cbb234, 32'hc24b179a} /* (7, 8, 24) {real, imag} */,
  {32'hc1e1171e, 32'h43187a20} /* (7, 8, 23) {real, imag} */,
  {32'h429d354a, 32'h4183eaa0} /* (7, 8, 22) {real, imag} */,
  {32'hc308d8ca, 32'hc255b398} /* (7, 8, 21) {real, imag} */,
  {32'hc287273b, 32'h41dd8efc} /* (7, 8, 20) {real, imag} */,
  {32'h41eeef6a, 32'hc1fd35e4} /* (7, 8, 19) {real, imag} */,
  {32'h42487d3e, 32'h41f1ed50} /* (7, 8, 18) {real, imag} */,
  {32'h41bc38a6, 32'h4238895c} /* (7, 8, 17) {real, imag} */,
  {32'h423e575c, 32'h00000000} /* (7, 8, 16) {real, imag} */,
  {32'h41bc38a6, 32'hc238895c} /* (7, 8, 15) {real, imag} */,
  {32'h42487d3e, 32'hc1f1ed50} /* (7, 8, 14) {real, imag} */,
  {32'h41eeef6a, 32'h41fd35e4} /* (7, 8, 13) {real, imag} */,
  {32'hc287273b, 32'hc1dd8efc} /* (7, 8, 12) {real, imag} */,
  {32'hc308d8ca, 32'h4255b398} /* (7, 8, 11) {real, imag} */,
  {32'h429d354a, 32'hc183eaa0} /* (7, 8, 10) {real, imag} */,
  {32'hc1e1171e, 32'hc3187a20} /* (7, 8, 9) {real, imag} */,
  {32'hc1cbb234, 32'h424b179a} /* (7, 8, 8) {real, imag} */,
  {32'h416702fa, 32'h4229cdbc} /* (7, 8, 7) {real, imag} */,
  {32'hc1aa397e, 32'hc29df706} /* (7, 8, 6) {real, imag} */,
  {32'hc33613fa, 32'hc3114998} /* (7, 8, 5) {real, imag} */,
  {32'h4330a681, 32'h4321128a} /* (7, 8, 4) {real, imag} */,
  {32'h434067a8, 32'hc30ff5c6} /* (7, 8, 3) {real, imag} */,
  {32'hc443b66b, 32'hc3e2279e} /* (7, 8, 2) {real, imag} */,
  {32'h450f6040, 32'h4485f3d4} /* (7, 8, 1) {real, imag} */,
  {32'h45251cf6, 32'h00000000} /* (7, 8, 0) {real, imag} */,
  {32'h452ace2f, 32'hc4a448a8} /* (7, 7, 31) {real, imag} */,
  {32'hc45eb0d8, 32'h4415bcda} /* (7, 7, 30) {real, imag} */,
  {32'h43522ad9, 32'hc1e46f64} /* (7, 7, 29) {real, imag} */,
  {32'h4327e850, 32'hc319646c} /* (7, 7, 28) {real, imag} */,
  {32'hc387944f, 32'h41d55cae} /* (7, 7, 27) {real, imag} */,
  {32'hc2d3748d, 32'hc1826621} /* (7, 7, 26) {real, imag} */,
  {32'h41a1568e, 32'hc31910fa} /* (7, 7, 25) {real, imag} */,
  {32'hc193eb8d, 32'hc1da1842} /* (7, 7, 24) {real, imag} */,
  {32'hc21c5d0b, 32'hc25323dc} /* (7, 7, 23) {real, imag} */,
  {32'hc193d93b, 32'h4288d5d0} /* (7, 7, 22) {real, imag} */,
  {32'hc23a1746, 32'h42e67e9f} /* (7, 7, 21) {real, imag} */,
  {32'h41a6e131, 32'h42515d20} /* (7, 7, 20) {real, imag} */,
  {32'h429f38b9, 32'h42255b6a} /* (7, 7, 19) {real, imag} */,
  {32'hc309b509, 32'h41f7b273} /* (7, 7, 18) {real, imag} */,
  {32'hc0a149e0, 32'hc0806778} /* (7, 7, 17) {real, imag} */,
  {32'h4223b238, 32'h00000000} /* (7, 7, 16) {real, imag} */,
  {32'hc0a149e0, 32'h40806778} /* (7, 7, 15) {real, imag} */,
  {32'hc309b509, 32'hc1f7b273} /* (7, 7, 14) {real, imag} */,
  {32'h429f38b9, 32'hc2255b6a} /* (7, 7, 13) {real, imag} */,
  {32'h41a6e131, 32'hc2515d20} /* (7, 7, 12) {real, imag} */,
  {32'hc23a1746, 32'hc2e67e9f} /* (7, 7, 11) {real, imag} */,
  {32'hc193d93b, 32'hc288d5d0} /* (7, 7, 10) {real, imag} */,
  {32'hc21c5d0b, 32'h425323dc} /* (7, 7, 9) {real, imag} */,
  {32'hc193eb8d, 32'h41da1842} /* (7, 7, 8) {real, imag} */,
  {32'h41a1568e, 32'h431910fa} /* (7, 7, 7) {real, imag} */,
  {32'hc2d3748d, 32'h41826621} /* (7, 7, 6) {real, imag} */,
  {32'hc387944f, 32'hc1d55cae} /* (7, 7, 5) {real, imag} */,
  {32'h4327e850, 32'h4319646c} /* (7, 7, 4) {real, imag} */,
  {32'h43522ad9, 32'h41e46f64} /* (7, 7, 3) {real, imag} */,
  {32'hc45eb0d8, 32'hc415bcda} /* (7, 7, 2) {real, imag} */,
  {32'h452ace2f, 32'h44a448a8} /* (7, 7, 1) {real, imag} */,
  {32'h4544dd04, 32'h00000000} /* (7, 7, 0) {real, imag} */,
  {32'h453b5b46, 32'hc4d8e070} /* (7, 6, 31) {real, imag} */,
  {32'hc427463a, 32'h442accd4} /* (7, 6, 30) {real, imag} */,
  {32'h426e7b9a, 32'h422a3c49} /* (7, 6, 29) {real, imag} */,
  {32'h430b6dd0, 32'hc1755c7c} /* (7, 6, 28) {real, imag} */,
  {32'hc323a93d, 32'h43000f8f} /* (7, 6, 27) {real, imag} */,
  {32'hc2810422, 32'h420d501c} /* (7, 6, 26) {real, imag} */,
  {32'h42b4e455, 32'hc309f206} /* (7, 6, 25) {real, imag} */,
  {32'hc2d70235, 32'h431de345} /* (7, 6, 24) {real, imag} */,
  {32'hc226c020, 32'h432a6504} /* (7, 6, 23) {real, imag} */,
  {32'hc30729be, 32'hc28ae391} /* (7, 6, 22) {real, imag} */,
  {32'hc2734d79, 32'h42a70938} /* (7, 6, 21) {real, imag} */,
  {32'h42c8eb9e, 32'hc0af78a4} /* (7, 6, 20) {real, imag} */,
  {32'h421bd222, 32'h420b7bf0} /* (7, 6, 19) {real, imag} */,
  {32'hc2a913e2, 32'h42a9fa87} /* (7, 6, 18) {real, imag} */,
  {32'hc1ffd13d, 32'hc26b25d2} /* (7, 6, 17) {real, imag} */,
  {32'h42d8db93, 32'h00000000} /* (7, 6, 16) {real, imag} */,
  {32'hc1ffd13d, 32'h426b25d2} /* (7, 6, 15) {real, imag} */,
  {32'hc2a913e2, 32'hc2a9fa87} /* (7, 6, 14) {real, imag} */,
  {32'h421bd222, 32'hc20b7bf0} /* (7, 6, 13) {real, imag} */,
  {32'h42c8eb9e, 32'h40af78a4} /* (7, 6, 12) {real, imag} */,
  {32'hc2734d79, 32'hc2a70938} /* (7, 6, 11) {real, imag} */,
  {32'hc30729be, 32'h428ae391} /* (7, 6, 10) {real, imag} */,
  {32'hc226c020, 32'hc32a6504} /* (7, 6, 9) {real, imag} */,
  {32'hc2d70235, 32'hc31de345} /* (7, 6, 8) {real, imag} */,
  {32'h42b4e455, 32'h4309f206} /* (7, 6, 7) {real, imag} */,
  {32'hc2810422, 32'hc20d501c} /* (7, 6, 6) {real, imag} */,
  {32'hc323a93d, 32'hc3000f8f} /* (7, 6, 5) {real, imag} */,
  {32'h430b6dd0, 32'h41755c7c} /* (7, 6, 4) {real, imag} */,
  {32'h426e7b9a, 32'hc22a3c49} /* (7, 6, 3) {real, imag} */,
  {32'hc427463a, 32'hc42accd4} /* (7, 6, 2) {real, imag} */,
  {32'h453b5b46, 32'h44d8e070} /* (7, 6, 1) {real, imag} */,
  {32'h456cdce6, 32'h00000000} /* (7, 6, 0) {real, imag} */,
  {32'h4531bf90, 32'hc5101f84} /* (7, 5, 31) {real, imag} */,
  {32'hc39f5ff6, 32'h4467f14d} /* (7, 5, 30) {real, imag} */,
  {32'h40e35324, 32'h41eafb1b} /* (7, 5, 29) {real, imag} */,
  {32'h413c38e8, 32'h436c70ea} /* (7, 5, 28) {real, imag} */,
  {32'hc33ef250, 32'h41c033c6} /* (7, 5, 27) {real, imag} */,
  {32'h42b75ee0, 32'h42ced9aa} /* (7, 5, 26) {real, imag} */,
  {32'h430204cc, 32'hc0b96390} /* (7, 5, 25) {real, imag} */,
  {32'h41428424, 32'h43005dce} /* (7, 5, 24) {real, imag} */,
  {32'hc27b44f3, 32'h42603d14} /* (7, 5, 23) {real, imag} */,
  {32'hc25c88b6, 32'h40336670} /* (7, 5, 22) {real, imag} */,
  {32'hc337a06c, 32'hc2142ad3} /* (7, 5, 21) {real, imag} */,
  {32'hc0ed1794, 32'hc130bfe8} /* (7, 5, 20) {real, imag} */,
  {32'hc256416d, 32'h40404340} /* (7, 5, 19) {real, imag} */,
  {32'hc2570efe, 32'hc2a1312e} /* (7, 5, 18) {real, imag} */,
  {32'hc185fd9d, 32'hc28723b0} /* (7, 5, 17) {real, imag} */,
  {32'hc28a443d, 32'h00000000} /* (7, 5, 16) {real, imag} */,
  {32'hc185fd9d, 32'h428723b0} /* (7, 5, 15) {real, imag} */,
  {32'hc2570efe, 32'h42a1312e} /* (7, 5, 14) {real, imag} */,
  {32'hc256416d, 32'hc0404340} /* (7, 5, 13) {real, imag} */,
  {32'hc0ed1794, 32'h4130bfe8} /* (7, 5, 12) {real, imag} */,
  {32'hc337a06c, 32'h42142ad3} /* (7, 5, 11) {real, imag} */,
  {32'hc25c88b6, 32'hc0336670} /* (7, 5, 10) {real, imag} */,
  {32'hc27b44f3, 32'hc2603d14} /* (7, 5, 9) {real, imag} */,
  {32'h41428424, 32'hc3005dce} /* (7, 5, 8) {real, imag} */,
  {32'h430204cc, 32'h40b96390} /* (7, 5, 7) {real, imag} */,
  {32'h42b75ee0, 32'hc2ced9aa} /* (7, 5, 6) {real, imag} */,
  {32'hc33ef250, 32'hc1c033c6} /* (7, 5, 5) {real, imag} */,
  {32'h413c38e8, 32'hc36c70ea} /* (7, 5, 4) {real, imag} */,
  {32'h40e35324, 32'hc1eafb1b} /* (7, 5, 3) {real, imag} */,
  {32'hc39f5ff6, 32'hc467f14d} /* (7, 5, 2) {real, imag} */,
  {32'h4531bf90, 32'h45101f84} /* (7, 5, 1) {real, imag} */,
  {32'h457d8496, 32'h00000000} /* (7, 5, 0) {real, imag} */,
  {32'h451caacd, 32'hc52bc1e5} /* (7, 4, 31) {real, imag} */,
  {32'h427e3898, 32'h44789206} /* (7, 4, 30) {real, imag} */,
  {32'h42661948, 32'hc21d02fa} /* (7, 4, 29) {real, imag} */,
  {32'h41fbf98c, 32'h436557c6} /* (7, 4, 28) {real, imag} */,
  {32'hc2dfb7d4, 32'hc1cd9a85} /* (7, 4, 27) {real, imag} */,
  {32'hc1c0f0ae, 32'h42e56e25} /* (7, 4, 26) {real, imag} */,
  {32'h42069f8e, 32'hc30aa1af} /* (7, 4, 25) {real, imag} */,
  {32'hc29095fe, 32'h41cbe277} /* (7, 4, 24) {real, imag} */,
  {32'hc1839185, 32'hc2a07816} /* (7, 4, 23) {real, imag} */,
  {32'h41efd774, 32'h42c55de5} /* (7, 4, 22) {real, imag} */,
  {32'hc1c6f3b2, 32'h42b0a12c} /* (7, 4, 21) {real, imag} */,
  {32'hc19e5294, 32'h4237d13b} /* (7, 4, 20) {real, imag} */,
  {32'hc1f4312a, 32'h42917c0b} /* (7, 4, 19) {real, imag} */,
  {32'h42ce7d43, 32'h42b9d9e2} /* (7, 4, 18) {real, imag} */,
  {32'hc1cd77c8, 32'h407bb850} /* (7, 4, 17) {real, imag} */,
  {32'hc259296c, 32'h00000000} /* (7, 4, 16) {real, imag} */,
  {32'hc1cd77c8, 32'hc07bb850} /* (7, 4, 15) {real, imag} */,
  {32'h42ce7d43, 32'hc2b9d9e2} /* (7, 4, 14) {real, imag} */,
  {32'hc1f4312a, 32'hc2917c0b} /* (7, 4, 13) {real, imag} */,
  {32'hc19e5294, 32'hc237d13b} /* (7, 4, 12) {real, imag} */,
  {32'hc1c6f3b2, 32'hc2b0a12c} /* (7, 4, 11) {real, imag} */,
  {32'h41efd774, 32'hc2c55de5} /* (7, 4, 10) {real, imag} */,
  {32'hc1839185, 32'h42a07816} /* (7, 4, 9) {real, imag} */,
  {32'hc29095fe, 32'hc1cbe277} /* (7, 4, 8) {real, imag} */,
  {32'h42069f8e, 32'h430aa1af} /* (7, 4, 7) {real, imag} */,
  {32'hc1c0f0ae, 32'hc2e56e25} /* (7, 4, 6) {real, imag} */,
  {32'hc2dfb7d4, 32'h41cd9a85} /* (7, 4, 5) {real, imag} */,
  {32'h41fbf98c, 32'hc36557c6} /* (7, 4, 4) {real, imag} */,
  {32'h42661948, 32'h421d02fa} /* (7, 4, 3) {real, imag} */,
  {32'h427e3898, 32'hc4789206} /* (7, 4, 2) {real, imag} */,
  {32'h451caacd, 32'h452bc1e5} /* (7, 4, 1) {real, imag} */,
  {32'h4588a70c, 32'h00000000} /* (7, 4, 0) {real, imag} */,
  {32'h4518a76c, 32'hc5386a85} /* (7, 3, 31) {real, imag} */,
  {32'h4396b5ea, 32'h44682ee4} /* (7, 3, 30) {real, imag} */,
  {32'h4233fb28, 32'h433ed196} /* (7, 3, 29) {real, imag} */,
  {32'hc29b4001, 32'h43b2ec00} /* (7, 3, 28) {real, imag} */,
  {32'hc35fa46d, 32'hc2bb76fd} /* (7, 3, 27) {real, imag} */,
  {32'hc24961bc, 32'hc2060d38} /* (7, 3, 26) {real, imag} */,
  {32'h3e7c1e00, 32'hc2c82882} /* (7, 3, 25) {real, imag} */,
  {32'hc20f2fd2, 32'h42258dfa} /* (7, 3, 24) {real, imag} */,
  {32'hc28edd9a, 32'hc202e7b0} /* (7, 3, 23) {real, imag} */,
  {32'hc2e740a8, 32'hc226f8a5} /* (7, 3, 22) {real, imag} */,
  {32'h42b38e71, 32'h41ed8afe} /* (7, 3, 21) {real, imag} */,
  {32'h42e630ea, 32'hc215d968} /* (7, 3, 20) {real, imag} */,
  {32'hc0ab5398, 32'h41cc5fcc} /* (7, 3, 19) {real, imag} */,
  {32'h41ff37e0, 32'h42979880} /* (7, 3, 18) {real, imag} */,
  {32'hc1ad162a, 32'h41829ea9} /* (7, 3, 17) {real, imag} */,
  {32'h42a8be9c, 32'h00000000} /* (7, 3, 16) {real, imag} */,
  {32'hc1ad162a, 32'hc1829ea9} /* (7, 3, 15) {real, imag} */,
  {32'h41ff37e0, 32'hc2979880} /* (7, 3, 14) {real, imag} */,
  {32'hc0ab5398, 32'hc1cc5fcc} /* (7, 3, 13) {real, imag} */,
  {32'h42e630ea, 32'h4215d968} /* (7, 3, 12) {real, imag} */,
  {32'h42b38e71, 32'hc1ed8afe} /* (7, 3, 11) {real, imag} */,
  {32'hc2e740a8, 32'h4226f8a5} /* (7, 3, 10) {real, imag} */,
  {32'hc28edd9a, 32'h4202e7b0} /* (7, 3, 9) {real, imag} */,
  {32'hc20f2fd2, 32'hc2258dfa} /* (7, 3, 8) {real, imag} */,
  {32'h3e7c1e00, 32'h42c82882} /* (7, 3, 7) {real, imag} */,
  {32'hc24961bc, 32'h42060d38} /* (7, 3, 6) {real, imag} */,
  {32'hc35fa46d, 32'h42bb76fd} /* (7, 3, 5) {real, imag} */,
  {32'hc29b4001, 32'hc3b2ec00} /* (7, 3, 4) {real, imag} */,
  {32'h4233fb28, 32'hc33ed196} /* (7, 3, 3) {real, imag} */,
  {32'h4396b5ea, 32'hc4682ee4} /* (7, 3, 2) {real, imag} */,
  {32'h4518a76c, 32'h45386a85} /* (7, 3, 1) {real, imag} */,
  {32'h458d17b5, 32'h00000000} /* (7, 3, 0) {real, imag} */,
  {32'h45133db4, 32'hc53d396b} /* (7, 2, 31) {real, imag} */,
  {32'h43c6cedf, 32'h445c5274} /* (7, 2, 30) {real, imag} */,
  {32'h4166ce38, 32'h42ed423a} /* (7, 2, 29) {real, imag} */,
  {32'hc3081f06, 32'h4393de68} /* (7, 2, 28) {real, imag} */,
  {32'hc31e5fe1, 32'hc1d29aa0} /* (7, 2, 27) {real, imag} */,
  {32'h41b5c24e, 32'hc26904ac} /* (7, 2, 26) {real, imag} */,
  {32'hc19a70d0, 32'hc258734f} /* (7, 2, 25) {real, imag} */,
  {32'h41cf0098, 32'h42f011be} /* (7, 2, 24) {real, imag} */,
  {32'h4281e300, 32'h428fb5e8} /* (7, 2, 23) {real, imag} */,
  {32'h41b478d5, 32'h4232f42d} /* (7, 2, 22) {real, imag} */,
  {32'hc0dac8f0, 32'h42362d2c} /* (7, 2, 21) {real, imag} */,
  {32'h40b5aaf4, 32'hc225ac0e} /* (7, 2, 20) {real, imag} */,
  {32'hc1a98e05, 32'hc0986130} /* (7, 2, 19) {real, imag} */,
  {32'hc1735eec, 32'hc044b824} /* (7, 2, 18) {real, imag} */,
  {32'h4193ec3e, 32'hc23c1fc0} /* (7, 2, 17) {real, imag} */,
  {32'h424137c0, 32'h00000000} /* (7, 2, 16) {real, imag} */,
  {32'h4193ec3e, 32'h423c1fc0} /* (7, 2, 15) {real, imag} */,
  {32'hc1735eec, 32'h4044b824} /* (7, 2, 14) {real, imag} */,
  {32'hc1a98e05, 32'h40986130} /* (7, 2, 13) {real, imag} */,
  {32'h40b5aaf4, 32'h4225ac0e} /* (7, 2, 12) {real, imag} */,
  {32'hc0dac8f0, 32'hc2362d2c} /* (7, 2, 11) {real, imag} */,
  {32'h41b478d5, 32'hc232f42d} /* (7, 2, 10) {real, imag} */,
  {32'h4281e300, 32'hc28fb5e8} /* (7, 2, 9) {real, imag} */,
  {32'h41cf0098, 32'hc2f011be} /* (7, 2, 8) {real, imag} */,
  {32'hc19a70d0, 32'h4258734f} /* (7, 2, 7) {real, imag} */,
  {32'h41b5c24e, 32'h426904ac} /* (7, 2, 6) {real, imag} */,
  {32'hc31e5fe1, 32'h41d29aa0} /* (7, 2, 5) {real, imag} */,
  {32'hc3081f06, 32'hc393de68} /* (7, 2, 4) {real, imag} */,
  {32'h4166ce38, 32'hc2ed423a} /* (7, 2, 3) {real, imag} */,
  {32'h43c6cedf, 32'hc45c5274} /* (7, 2, 2) {real, imag} */,
  {32'h45133db4, 32'h453d396b} /* (7, 2, 1) {real, imag} */,
  {32'h459434b6, 32'h00000000} /* (7, 2, 0) {real, imag} */,
  {32'h45154b8e, 32'hc52ee45c} /* (7, 1, 31) {real, imag} */,
  {32'h43b56681, 32'h4443c58a} /* (7, 1, 30) {real, imag} */,
  {32'hc32cd73e, 32'h428cab81} /* (7, 1, 29) {real, imag} */,
  {32'hc2cca31b, 32'h43388af0} /* (7, 1, 28) {real, imag} */,
  {32'hc28079a1, 32'h4196f4fa} /* (7, 1, 27) {real, imag} */,
  {32'hc2e7b6f2, 32'h424a9bb1} /* (7, 1, 26) {real, imag} */,
  {32'hc1937076, 32'hc2913bc8} /* (7, 1, 25) {real, imag} */,
  {32'h42595d16, 32'h429da270} /* (7, 1, 24) {real, imag} */,
  {32'h42a7a8bb, 32'hc2c922b6} /* (7, 1, 23) {real, imag} */,
  {32'h42798ebe, 32'h41dfe301} /* (7, 1, 22) {real, imag} */,
  {32'h4261867c, 32'h4304374f} /* (7, 1, 21) {real, imag} */,
  {32'hc2920d88, 32'h4214743c} /* (7, 1, 20) {real, imag} */,
  {32'hc2896140, 32'h4271a35a} /* (7, 1, 19) {real, imag} */,
  {32'h42a5bc08, 32'h41aed796} /* (7, 1, 18) {real, imag} */,
  {32'hc1cc8bb6, 32'hc1843b46} /* (7, 1, 17) {real, imag} */,
  {32'h3f883a40, 32'h00000000} /* (7, 1, 16) {real, imag} */,
  {32'hc1cc8bb6, 32'h41843b46} /* (7, 1, 15) {real, imag} */,
  {32'h42a5bc08, 32'hc1aed796} /* (7, 1, 14) {real, imag} */,
  {32'hc2896140, 32'hc271a35a} /* (7, 1, 13) {real, imag} */,
  {32'hc2920d88, 32'hc214743c} /* (7, 1, 12) {real, imag} */,
  {32'h4261867c, 32'hc304374f} /* (7, 1, 11) {real, imag} */,
  {32'h42798ebe, 32'hc1dfe301} /* (7, 1, 10) {real, imag} */,
  {32'h42a7a8bb, 32'h42c922b6} /* (7, 1, 9) {real, imag} */,
  {32'h42595d16, 32'hc29da270} /* (7, 1, 8) {real, imag} */,
  {32'hc1937076, 32'h42913bc8} /* (7, 1, 7) {real, imag} */,
  {32'hc2e7b6f2, 32'hc24a9bb1} /* (7, 1, 6) {real, imag} */,
  {32'hc28079a1, 32'hc196f4fa} /* (7, 1, 5) {real, imag} */,
  {32'hc2cca31b, 32'hc3388af0} /* (7, 1, 4) {real, imag} */,
  {32'hc32cd73e, 32'hc28cab81} /* (7, 1, 3) {real, imag} */,
  {32'h43b56681, 32'hc443c58a} /* (7, 1, 2) {real, imag} */,
  {32'h45154b8e, 32'h452ee45c} /* (7, 1, 1) {real, imag} */,
  {32'h4591cf8c, 32'h00000000} /* (7, 1, 0) {real, imag} */,
  {32'h4521c640, 32'hc50853a3} /* (7, 0, 31) {real, imag} */,
  {32'h4152cc00, 32'h441aec3c} /* (7, 0, 30) {real, imag} */,
  {32'hc311e958, 32'hc2903db2} /* (7, 0, 29) {real, imag} */,
  {32'h41411650, 32'h431d1a94} /* (7, 0, 28) {real, imag} */,
  {32'hc07d2590, 32'hc0e0b57c} /* (7, 0, 27) {real, imag} */,
  {32'h4189cc67, 32'hc1d15864} /* (7, 0, 26) {real, imag} */,
  {32'hc2326228, 32'hc245f4a4} /* (7, 0, 25) {real, imag} */,
  {32'hc29e2388, 32'hc241cefc} /* (7, 0, 24) {real, imag} */,
  {32'hc1d44d30, 32'hc277891d} /* (7, 0, 23) {real, imag} */,
  {32'h425d487e, 32'hc15965b0} /* (7, 0, 22) {real, imag} */,
  {32'h41cbb25e, 32'hc1c87834} /* (7, 0, 21) {real, imag} */,
  {32'h41e7edce, 32'hc0739290} /* (7, 0, 20) {real, imag} */,
  {32'h41c511ca, 32'h42d96f08} /* (7, 0, 19) {real, imag} */,
  {32'hc2bde81b, 32'hc1245c25} /* (7, 0, 18) {real, imag} */,
  {32'hbff9cb68, 32'hc10c02b4} /* (7, 0, 17) {real, imag} */,
  {32'hc0e95fa8, 32'h00000000} /* (7, 0, 16) {real, imag} */,
  {32'hbff9cb68, 32'h410c02b4} /* (7, 0, 15) {real, imag} */,
  {32'hc2bde81b, 32'h41245c25} /* (7, 0, 14) {real, imag} */,
  {32'h41c511ca, 32'hc2d96f08} /* (7, 0, 13) {real, imag} */,
  {32'h41e7edce, 32'h40739290} /* (7, 0, 12) {real, imag} */,
  {32'h41cbb25e, 32'h41c87834} /* (7, 0, 11) {real, imag} */,
  {32'h425d487e, 32'h415965b0} /* (7, 0, 10) {real, imag} */,
  {32'hc1d44d30, 32'h4277891d} /* (7, 0, 9) {real, imag} */,
  {32'hc29e2388, 32'h4241cefc} /* (7, 0, 8) {real, imag} */,
  {32'hc2326228, 32'h4245f4a4} /* (7, 0, 7) {real, imag} */,
  {32'h4189cc67, 32'h41d15864} /* (7, 0, 6) {real, imag} */,
  {32'hc07d2590, 32'h40e0b57c} /* (7, 0, 5) {real, imag} */,
  {32'h41411650, 32'hc31d1a94} /* (7, 0, 4) {real, imag} */,
  {32'hc311e958, 32'h42903db2} /* (7, 0, 3) {real, imag} */,
  {32'h4152cc00, 32'hc41aec3c} /* (7, 0, 2) {real, imag} */,
  {32'h4521c640, 32'h450853a3} /* (7, 0, 1) {real, imag} */,
  {32'h4587a5ea, 32'h00000000} /* (7, 0, 0) {real, imag} */,
  {32'h4507a6e6, 32'hc48fed82} /* (6, 31, 31) {real, imag} */,
  {32'hc386a740, 32'h431164a8} /* (6, 31, 30) {real, imag} */,
  {32'h42001704, 32'h416c2b28} /* (6, 31, 29) {real, imag} */,
  {32'h42b85e80, 32'h421a0173} /* (6, 31, 28) {real, imag} */,
  {32'hc2560a4d, 32'h40bf46fc} /* (6, 31, 27) {real, imag} */,
  {32'hc1693588, 32'hc10d4ede} /* (6, 31, 26) {real, imag} */,
  {32'h41ed11ed, 32'h416412f4} /* (6, 31, 25) {real, imag} */,
  {32'h40e527cc, 32'h4257d07e} /* (6, 31, 24) {real, imag} */,
  {32'h4205cea3, 32'hc1708582} /* (6, 31, 23) {real, imag} */,
  {32'h419220aa, 32'hc200c528} /* (6, 31, 22) {real, imag} */,
  {32'h419b7db9, 32'h41da3f03} /* (6, 31, 21) {real, imag} */,
  {32'hc10faa60, 32'h40d52054} /* (6, 31, 20) {real, imag} */,
  {32'h420251b2, 32'h42d0e25c} /* (6, 31, 19) {real, imag} */,
  {32'hc1d4102d, 32'h429ff183} /* (6, 31, 18) {real, imag} */,
  {32'h420795f0, 32'hc04c6eda} /* (6, 31, 17) {real, imag} */,
  {32'h42225610, 32'h00000000} /* (6, 31, 16) {real, imag} */,
  {32'h420795f0, 32'h404c6eda} /* (6, 31, 15) {real, imag} */,
  {32'hc1d4102d, 32'hc29ff183} /* (6, 31, 14) {real, imag} */,
  {32'h420251b2, 32'hc2d0e25c} /* (6, 31, 13) {real, imag} */,
  {32'hc10faa60, 32'hc0d52054} /* (6, 31, 12) {real, imag} */,
  {32'h419b7db9, 32'hc1da3f03} /* (6, 31, 11) {real, imag} */,
  {32'h419220aa, 32'h4200c528} /* (6, 31, 10) {real, imag} */,
  {32'h4205cea3, 32'h41708582} /* (6, 31, 9) {real, imag} */,
  {32'h40e527cc, 32'hc257d07e} /* (6, 31, 8) {real, imag} */,
  {32'h41ed11ed, 32'hc16412f4} /* (6, 31, 7) {real, imag} */,
  {32'hc1693588, 32'h410d4ede} /* (6, 31, 6) {real, imag} */,
  {32'hc2560a4d, 32'hc0bf46fc} /* (6, 31, 5) {real, imag} */,
  {32'h42b85e80, 32'hc21a0173} /* (6, 31, 4) {real, imag} */,
  {32'h42001704, 32'hc16c2b28} /* (6, 31, 3) {real, imag} */,
  {32'hc386a740, 32'hc31164a8} /* (6, 31, 2) {real, imag} */,
  {32'h4507a6e6, 32'h448fed82} /* (6, 31, 1) {real, imag} */,
  {32'h4557527f, 32'h00000000} /* (6, 31, 0) {real, imag} */,
  {32'h45295e30, 32'hc476467d} /* (6, 30, 31) {real, imag} */,
  {32'hc3ec2662, 32'h43088662} /* (6, 30, 30) {real, imag} */,
  {32'h42a4aab3, 32'h400843a0} /* (6, 30, 29) {real, imag} */,
  {32'h42c68b46, 32'hbe491b00} /* (6, 30, 28) {real, imag} */,
  {32'hc35c9ccc, 32'hc236eb61} /* (6, 30, 27) {real, imag} */,
  {32'h418dbdac, 32'h42f91df3} /* (6, 30, 26) {real, imag} */,
  {32'hc2998ecc, 32'hc2517a26} /* (6, 30, 25) {real, imag} */,
  {32'hc2a1e0fb, 32'h41d9127c} /* (6, 30, 24) {real, imag} */,
  {32'hc18b5eca, 32'h42b45621} /* (6, 30, 23) {real, imag} */,
  {32'h42aee690, 32'hc2b6ca9d} /* (6, 30, 22) {real, imag} */,
  {32'hc2f0cad9, 32'h430919b8} /* (6, 30, 21) {real, imag} */,
  {32'h41e25432, 32'hc284478e} /* (6, 30, 20) {real, imag} */,
  {32'h4250a25b, 32'h42211fc4} /* (6, 30, 19) {real, imag} */,
  {32'hc2802adb, 32'h42328ec9} /* (6, 30, 18) {real, imag} */,
  {32'h414d827c, 32'h422d7af1} /* (6, 30, 17) {real, imag} */,
  {32'hc0f05aa4, 32'h00000000} /* (6, 30, 16) {real, imag} */,
  {32'h414d827c, 32'hc22d7af1} /* (6, 30, 15) {real, imag} */,
  {32'hc2802adb, 32'hc2328ec9} /* (6, 30, 14) {real, imag} */,
  {32'h4250a25b, 32'hc2211fc4} /* (6, 30, 13) {real, imag} */,
  {32'h41e25432, 32'h4284478e} /* (6, 30, 12) {real, imag} */,
  {32'hc2f0cad9, 32'hc30919b8} /* (6, 30, 11) {real, imag} */,
  {32'h42aee690, 32'h42b6ca9d} /* (6, 30, 10) {real, imag} */,
  {32'hc18b5eca, 32'hc2b45621} /* (6, 30, 9) {real, imag} */,
  {32'hc2a1e0fb, 32'hc1d9127c} /* (6, 30, 8) {real, imag} */,
  {32'hc2998ecc, 32'h42517a26} /* (6, 30, 7) {real, imag} */,
  {32'h418dbdac, 32'hc2f91df3} /* (6, 30, 6) {real, imag} */,
  {32'hc35c9ccc, 32'h4236eb61} /* (6, 30, 5) {real, imag} */,
  {32'h42c68b46, 32'h3e491b00} /* (6, 30, 4) {real, imag} */,
  {32'h42a4aab3, 32'hc00843a0} /* (6, 30, 3) {real, imag} */,
  {32'hc3ec2662, 32'hc3088662} /* (6, 30, 2) {real, imag} */,
  {32'h45295e30, 32'h4476467d} /* (6, 30, 1) {real, imag} */,
  {32'h45598b5d, 32'h00000000} /* (6, 30, 0) {real, imag} */,
  {32'h451e9cf1, 32'hc41abd58} /* (6, 29, 31) {real, imag} */,
  {32'hc423c16e, 32'h43568192} /* (6, 29, 30) {real, imag} */,
  {32'h4291ece8, 32'hc32beecb} /* (6, 29, 29) {real, imag} */,
  {32'h431d2241, 32'hc31d2b62} /* (6, 29, 28) {real, imag} */,
  {32'hc32ead86, 32'h42536a97} /* (6, 29, 27) {real, imag} */,
  {32'h42580b5f, 32'h41cefed1} /* (6, 29, 26) {real, imag} */,
  {32'h422f233e, 32'hc224b671} /* (6, 29, 25) {real, imag} */,
  {32'h41c3718c, 32'h41dc216b} /* (6, 29, 24) {real, imag} */,
  {32'hc2321a4c, 32'h42afc5bc} /* (6, 29, 23) {real, imag} */,
  {32'hc1de2b13, 32'h417bccf2} /* (6, 29, 22) {real, imag} */,
  {32'hc09410f8, 32'h42b1cfdd} /* (6, 29, 21) {real, imag} */,
  {32'hc1a3ef76, 32'h40a24c14} /* (6, 29, 20) {real, imag} */,
  {32'hc28c93f6, 32'hc24a31d4} /* (6, 29, 19) {real, imag} */,
  {32'hc2976432, 32'h4245b8d1} /* (6, 29, 18) {real, imag} */,
  {32'h41ba205e, 32'hc19299dc} /* (6, 29, 17) {real, imag} */,
  {32'h422ea4b2, 32'h00000000} /* (6, 29, 16) {real, imag} */,
  {32'h41ba205e, 32'h419299dc} /* (6, 29, 15) {real, imag} */,
  {32'hc2976432, 32'hc245b8d1} /* (6, 29, 14) {real, imag} */,
  {32'hc28c93f6, 32'h424a31d4} /* (6, 29, 13) {real, imag} */,
  {32'hc1a3ef76, 32'hc0a24c14} /* (6, 29, 12) {real, imag} */,
  {32'hc09410f8, 32'hc2b1cfdd} /* (6, 29, 11) {real, imag} */,
  {32'hc1de2b13, 32'hc17bccf2} /* (6, 29, 10) {real, imag} */,
  {32'hc2321a4c, 32'hc2afc5bc} /* (6, 29, 9) {real, imag} */,
  {32'h41c3718c, 32'hc1dc216b} /* (6, 29, 8) {real, imag} */,
  {32'h422f233e, 32'h4224b671} /* (6, 29, 7) {real, imag} */,
  {32'h42580b5f, 32'hc1cefed1} /* (6, 29, 6) {real, imag} */,
  {32'hc32ead86, 32'hc2536a97} /* (6, 29, 5) {real, imag} */,
  {32'h431d2241, 32'h431d2b62} /* (6, 29, 4) {real, imag} */,
  {32'h4291ece8, 32'h432beecb} /* (6, 29, 3) {real, imag} */,
  {32'hc423c16e, 32'hc3568192} /* (6, 29, 2) {real, imag} */,
  {32'h451e9cf1, 32'h441abd58} /* (6, 29, 1) {real, imag} */,
  {32'h456062f0, 32'h00000000} /* (6, 29, 0) {real, imag} */,
  {32'h451eac1b, 32'hc3b0abd8} /* (6, 28, 31) {real, imag} */,
  {32'hc44a4f73, 32'h43945340} /* (6, 28, 30) {real, imag} */,
  {32'h4298c8d9, 32'hc2482dee} /* (6, 28, 29) {real, imag} */,
  {32'h42c8e183, 32'hc292c458} /* (6, 28, 28) {real, imag} */,
  {32'hc3a14ad2, 32'h42840d9c} /* (6, 28, 27) {real, imag} */,
  {32'hc1a9018e, 32'hc1d428a0} /* (6, 28, 26) {real, imag} */,
  {32'h421fe9e1, 32'hc27fe680} /* (6, 28, 25) {real, imag} */,
  {32'hc1a4982d, 32'h41a71362} /* (6, 28, 24) {real, imag} */,
  {32'hc26e63f0, 32'hc223232c} /* (6, 28, 23) {real, imag} */,
  {32'h41b98a2a, 32'hc28ac41b} /* (6, 28, 22) {real, imag} */,
  {32'hc1f3cf87, 32'h42cb9d6a} /* (6, 28, 21) {real, imag} */,
  {32'h42a71ce8, 32'hc24c8e66} /* (6, 28, 20) {real, imag} */,
  {32'h41d3e400, 32'hc1185e2c} /* (6, 28, 19) {real, imag} */,
  {32'h4131d91b, 32'h42b5e0b9} /* (6, 28, 18) {real, imag} */,
  {32'h40d9fa38, 32'hc2017ea6} /* (6, 28, 17) {real, imag} */,
  {32'hc1a25595, 32'h00000000} /* (6, 28, 16) {real, imag} */,
  {32'h40d9fa38, 32'h42017ea6} /* (6, 28, 15) {real, imag} */,
  {32'h4131d91b, 32'hc2b5e0b9} /* (6, 28, 14) {real, imag} */,
  {32'h41d3e400, 32'h41185e2c} /* (6, 28, 13) {real, imag} */,
  {32'h42a71ce8, 32'h424c8e66} /* (6, 28, 12) {real, imag} */,
  {32'hc1f3cf87, 32'hc2cb9d6a} /* (6, 28, 11) {real, imag} */,
  {32'h41b98a2a, 32'h428ac41b} /* (6, 28, 10) {real, imag} */,
  {32'hc26e63f0, 32'h4223232c} /* (6, 28, 9) {real, imag} */,
  {32'hc1a4982d, 32'hc1a71362} /* (6, 28, 8) {real, imag} */,
  {32'h421fe9e1, 32'h427fe680} /* (6, 28, 7) {real, imag} */,
  {32'hc1a9018e, 32'h41d428a0} /* (6, 28, 6) {real, imag} */,
  {32'hc3a14ad2, 32'hc2840d9c} /* (6, 28, 5) {real, imag} */,
  {32'h42c8e183, 32'h4292c458} /* (6, 28, 4) {real, imag} */,
  {32'h4298c8d9, 32'h42482dee} /* (6, 28, 3) {real, imag} */,
  {32'hc44a4f73, 32'hc3945340} /* (6, 28, 2) {real, imag} */,
  {32'h451eac1b, 32'h43b0abd8} /* (6, 28, 1) {real, imag} */,
  {32'h455c4b3a, 32'h00000000} /* (6, 28, 0) {real, imag} */,
  {32'h451c98cc, 32'hc3deda76} /* (6, 27, 31) {real, imag} */,
  {32'hc457b72d, 32'h43964a55} /* (6, 27, 30) {real, imag} */,
  {32'h42956521, 32'h420fd121} /* (6, 27, 29) {real, imag} */,
  {32'h431fae8e, 32'hc32f11cd} /* (6, 27, 28) {real, imag} */,
  {32'hc351da10, 32'h424ab146} /* (6, 27, 27) {real, imag} */,
  {32'h42b63638, 32'h4247e9ca} /* (6, 27, 26) {real, imag} */,
  {32'h413136e8, 32'h40eeb6a0} /* (6, 27, 25) {real, imag} */,
  {32'hc2570b66, 32'hc20d2c24} /* (6, 27, 24) {real, imag} */,
  {32'h42341264, 32'hc13b7c1c} /* (6, 27, 23) {real, imag} */,
  {32'hc21fa8bc, 32'h41aebeaa} /* (6, 27, 22) {real, imag} */,
  {32'hc1f7b278, 32'h40de8634} /* (6, 27, 21) {real, imag} */,
  {32'h428a3ad4, 32'hbfb11ab8} /* (6, 27, 20) {real, imag} */,
  {32'h42278daa, 32'hc1ee31b9} /* (6, 27, 19) {real, imag} */,
  {32'hc2bac404, 32'h42f68ff2} /* (6, 27, 18) {real, imag} */,
  {32'hbf3776c0, 32'hc1ce3278} /* (6, 27, 17) {real, imag} */,
  {32'h421ac9e2, 32'h00000000} /* (6, 27, 16) {real, imag} */,
  {32'hbf3776c0, 32'h41ce3278} /* (6, 27, 15) {real, imag} */,
  {32'hc2bac404, 32'hc2f68ff2} /* (6, 27, 14) {real, imag} */,
  {32'h42278daa, 32'h41ee31b9} /* (6, 27, 13) {real, imag} */,
  {32'h428a3ad4, 32'h3fb11ab8} /* (6, 27, 12) {real, imag} */,
  {32'hc1f7b278, 32'hc0de8634} /* (6, 27, 11) {real, imag} */,
  {32'hc21fa8bc, 32'hc1aebeaa} /* (6, 27, 10) {real, imag} */,
  {32'h42341264, 32'h413b7c1c} /* (6, 27, 9) {real, imag} */,
  {32'hc2570b66, 32'h420d2c24} /* (6, 27, 8) {real, imag} */,
  {32'h413136e8, 32'hc0eeb6a0} /* (6, 27, 7) {real, imag} */,
  {32'h42b63638, 32'hc247e9ca} /* (6, 27, 6) {real, imag} */,
  {32'hc351da10, 32'hc24ab146} /* (6, 27, 5) {real, imag} */,
  {32'h431fae8e, 32'h432f11cd} /* (6, 27, 4) {real, imag} */,
  {32'h42956521, 32'hc20fd121} /* (6, 27, 3) {real, imag} */,
  {32'hc457b72d, 32'hc3964a55} /* (6, 27, 2) {real, imag} */,
  {32'h451c98cc, 32'h43deda76} /* (6, 27, 1) {real, imag} */,
  {32'h454fb75b, 32'h00000000} /* (6, 27, 0) {real, imag} */,
  {32'h45130850, 32'hc394ad76} /* (6, 26, 31) {real, imag} */,
  {32'hc45be24a, 32'h4313e0a5} /* (6, 26, 30) {real, imag} */,
  {32'hc18775c4, 32'hc30f3216} /* (6, 26, 29) {real, imag} */,
  {32'h42ffeb5f, 32'hc2d07310} /* (6, 26, 28) {real, imag} */,
  {32'hc33dee41, 32'h42f23e8b} /* (6, 26, 27) {real, imag} */,
  {32'h42fc02bb, 32'hc23ce964} /* (6, 26, 26) {real, imag} */,
  {32'h41cdb46c, 32'h41f4a6b6} /* (6, 26, 25) {real, imag} */,
  {32'hbe675700, 32'h42932393} /* (6, 26, 24) {real, imag} */,
  {32'hc19b6c2a, 32'h429d693a} /* (6, 26, 23) {real, imag} */,
  {32'h416f4852, 32'hc22c7cba} /* (6, 26, 22) {real, imag} */,
  {32'h40be7c10, 32'h42536000} /* (6, 26, 21) {real, imag} */,
  {32'hc214c0b8, 32'hc1e07dce} /* (6, 26, 20) {real, imag} */,
  {32'hc17b55ae, 32'hc2c1c18c} /* (6, 26, 19) {real, imag} */,
  {32'hc23541d3, 32'h425e4f2c} /* (6, 26, 18) {real, imag} */,
  {32'hc26312ce, 32'hc19f73a8} /* (6, 26, 17) {real, imag} */,
  {32'hc11f38cd, 32'h00000000} /* (6, 26, 16) {real, imag} */,
  {32'hc26312ce, 32'h419f73a8} /* (6, 26, 15) {real, imag} */,
  {32'hc23541d3, 32'hc25e4f2c} /* (6, 26, 14) {real, imag} */,
  {32'hc17b55ae, 32'h42c1c18c} /* (6, 26, 13) {real, imag} */,
  {32'hc214c0b8, 32'h41e07dce} /* (6, 26, 12) {real, imag} */,
  {32'h40be7c10, 32'hc2536000} /* (6, 26, 11) {real, imag} */,
  {32'h416f4852, 32'h422c7cba} /* (6, 26, 10) {real, imag} */,
  {32'hc19b6c2a, 32'hc29d693a} /* (6, 26, 9) {real, imag} */,
  {32'hbe675700, 32'hc2932393} /* (6, 26, 8) {real, imag} */,
  {32'h41cdb46c, 32'hc1f4a6b6} /* (6, 26, 7) {real, imag} */,
  {32'h42fc02bb, 32'h423ce964} /* (6, 26, 6) {real, imag} */,
  {32'hc33dee41, 32'hc2f23e8b} /* (6, 26, 5) {real, imag} */,
  {32'h42ffeb5f, 32'h42d07310} /* (6, 26, 4) {real, imag} */,
  {32'hc18775c4, 32'h430f3216} /* (6, 26, 3) {real, imag} */,
  {32'hc45be24a, 32'hc313e0a5} /* (6, 26, 2) {real, imag} */,
  {32'h45130850, 32'h4394ad76} /* (6, 26, 1) {real, imag} */,
  {32'h453f8da8, 32'h00000000} /* (6, 26, 0) {real, imag} */,
  {32'h4508a9c1, 32'hc391dd51} /* (6, 25, 31) {real, imag} */,
  {32'hc44e24e9, 32'h4307fecb} /* (6, 25, 30) {real, imag} */,
  {32'h4256c334, 32'hc2bf78e6} /* (6, 25, 29) {real, imag} */,
  {32'h42955817, 32'hc1846be6} /* (6, 25, 28) {real, imag} */,
  {32'hc2a90ea2, 32'h42b3923a} /* (6, 25, 27) {real, imag} */,
  {32'h4243d390, 32'hc30e3216} /* (6, 25, 26) {real, imag} */,
  {32'hc0c84e6a, 32'h421d610f} /* (6, 25, 25) {real, imag} */,
  {32'hc321f48a, 32'h42838bce} /* (6, 25, 24) {real, imag} */,
  {32'hc2a78e64, 32'h41e0aa84} /* (6, 25, 23) {real, imag} */,
  {32'h4197e22e, 32'h40925e58} /* (6, 25, 22) {real, imag} */,
  {32'hc29ce3d1, 32'h42153494} /* (6, 25, 21) {real, imag} */,
  {32'h42125ea4, 32'hc1b9c8ea} /* (6, 25, 20) {real, imag} */,
  {32'hc2a8c309, 32'hc139d3e2} /* (6, 25, 19) {real, imag} */,
  {32'h42082859, 32'h4271c919} /* (6, 25, 18) {real, imag} */,
  {32'hc16fc424, 32'h429bf61c} /* (6, 25, 17) {real, imag} */,
  {32'hc1164408, 32'h00000000} /* (6, 25, 16) {real, imag} */,
  {32'hc16fc424, 32'hc29bf61c} /* (6, 25, 15) {real, imag} */,
  {32'h42082859, 32'hc271c919} /* (6, 25, 14) {real, imag} */,
  {32'hc2a8c309, 32'h4139d3e2} /* (6, 25, 13) {real, imag} */,
  {32'h42125ea4, 32'h41b9c8ea} /* (6, 25, 12) {real, imag} */,
  {32'hc29ce3d1, 32'hc2153494} /* (6, 25, 11) {real, imag} */,
  {32'h4197e22e, 32'hc0925e58} /* (6, 25, 10) {real, imag} */,
  {32'hc2a78e64, 32'hc1e0aa84} /* (6, 25, 9) {real, imag} */,
  {32'hc321f48a, 32'hc2838bce} /* (6, 25, 8) {real, imag} */,
  {32'hc0c84e6a, 32'hc21d610f} /* (6, 25, 7) {real, imag} */,
  {32'h4243d390, 32'h430e3216} /* (6, 25, 6) {real, imag} */,
  {32'hc2a90ea2, 32'hc2b3923a} /* (6, 25, 5) {real, imag} */,
  {32'h42955817, 32'h41846be6} /* (6, 25, 4) {real, imag} */,
  {32'h4256c334, 32'h42bf78e6} /* (6, 25, 3) {real, imag} */,
  {32'hc44e24e9, 32'hc307fecb} /* (6, 25, 2) {real, imag} */,
  {32'h4508a9c1, 32'h4391dd51} /* (6, 25, 1) {real, imag} */,
  {32'h4532e6f2, 32'h00000000} /* (6, 25, 0) {real, imag} */,
  {32'h44eb9357, 32'hc398fd54} /* (6, 24, 31) {real, imag} */,
  {32'hc43f40c5, 32'h4301d44c} /* (6, 24, 30) {real, imag} */,
  {32'h41a99b68, 32'hc21434b1} /* (6, 24, 29) {real, imag} */,
  {32'h3ff62340, 32'hc2030883} /* (6, 24, 28) {real, imag} */,
  {32'hc2db7584, 32'h42493860} /* (6, 24, 27) {real, imag} */,
  {32'hc0e49d90, 32'hc215fccc} /* (6, 24, 26) {real, imag} */,
  {32'h42bce716, 32'h4129a5c0} /* (6, 24, 25) {real, imag} */,
  {32'hc2b1db51, 32'h427558a2} /* (6, 24, 24) {real, imag} */,
  {32'hc18fcd6d, 32'hc1dfb8ec} /* (6, 24, 23) {real, imag} */,
  {32'hc2c756ca, 32'hc14c0efa} /* (6, 24, 22) {real, imag} */,
  {32'hc1c8324e, 32'h427548b2} /* (6, 24, 21) {real, imag} */,
  {32'h424857b6, 32'hc31f4774} /* (6, 24, 20) {real, imag} */,
  {32'h42af3eb6, 32'h42b9317a} /* (6, 24, 19) {real, imag} */,
  {32'h41e7a0a7, 32'h423d1ba7} /* (6, 24, 18) {real, imag} */,
  {32'h41869b98, 32'hc0f7f894} /* (6, 24, 17) {real, imag} */,
  {32'h4205c26f, 32'h00000000} /* (6, 24, 16) {real, imag} */,
  {32'h41869b98, 32'h40f7f894} /* (6, 24, 15) {real, imag} */,
  {32'h41e7a0a7, 32'hc23d1ba7} /* (6, 24, 14) {real, imag} */,
  {32'h42af3eb6, 32'hc2b9317a} /* (6, 24, 13) {real, imag} */,
  {32'h424857b6, 32'h431f4774} /* (6, 24, 12) {real, imag} */,
  {32'hc1c8324e, 32'hc27548b2} /* (6, 24, 11) {real, imag} */,
  {32'hc2c756ca, 32'h414c0efa} /* (6, 24, 10) {real, imag} */,
  {32'hc18fcd6d, 32'h41dfb8ec} /* (6, 24, 9) {real, imag} */,
  {32'hc2b1db51, 32'hc27558a2} /* (6, 24, 8) {real, imag} */,
  {32'h42bce716, 32'hc129a5c0} /* (6, 24, 7) {real, imag} */,
  {32'hc0e49d90, 32'h4215fccc} /* (6, 24, 6) {real, imag} */,
  {32'hc2db7584, 32'hc2493860} /* (6, 24, 5) {real, imag} */,
  {32'h3ff62340, 32'h42030883} /* (6, 24, 4) {real, imag} */,
  {32'h41a99b68, 32'h421434b1} /* (6, 24, 3) {real, imag} */,
  {32'hc43f40c5, 32'hc301d44c} /* (6, 24, 2) {real, imag} */,
  {32'h44eb9357, 32'h4398fd54} /* (6, 24, 1) {real, imag} */,
  {32'h4526973a, 32'h00000000} /* (6, 24, 0) {real, imag} */,
  {32'h44afb9df, 32'hc3cad4d7} /* (6, 23, 31) {real, imag} */,
  {32'hc4236a69, 32'h42808a6a} /* (6, 23, 30) {real, imag} */,
  {32'h4229cce3, 32'hc2eb0f83} /* (6, 23, 29) {real, imag} */,
  {32'h426166c0, 32'hc22a60d8} /* (6, 23, 28) {real, imag} */,
  {32'hc2861237, 32'h40552a80} /* (6, 23, 27) {real, imag} */,
  {32'hc1858e1b, 32'hc2a6bbd3} /* (6, 23, 26) {real, imag} */,
  {32'hc1b0a85e, 32'hc275a488} /* (6, 23, 25) {real, imag} */,
  {32'hc2947597, 32'hc24f47ac} /* (6, 23, 24) {real, imag} */,
  {32'h41a6671f, 32'h42ac1d82} /* (6, 23, 23) {real, imag} */,
  {32'hc28a109c, 32'h40e8103c} /* (6, 23, 22) {real, imag} */,
  {32'hc17e0140, 32'h425c7e48} /* (6, 23, 21) {real, imag} */,
  {32'h4071cba8, 32'hc209665e} /* (6, 23, 20) {real, imag} */,
  {32'h41e03829, 32'h42436d68} /* (6, 23, 19) {real, imag} */,
  {32'hc26b5fc3, 32'hc25f12bc} /* (6, 23, 18) {real, imag} */,
  {32'h41ffc7a4, 32'hc213352c} /* (6, 23, 17) {real, imag} */,
  {32'h41890fde, 32'h00000000} /* (6, 23, 16) {real, imag} */,
  {32'h41ffc7a4, 32'h4213352c} /* (6, 23, 15) {real, imag} */,
  {32'hc26b5fc3, 32'h425f12bc} /* (6, 23, 14) {real, imag} */,
  {32'h41e03829, 32'hc2436d68} /* (6, 23, 13) {real, imag} */,
  {32'h4071cba8, 32'h4209665e} /* (6, 23, 12) {real, imag} */,
  {32'hc17e0140, 32'hc25c7e48} /* (6, 23, 11) {real, imag} */,
  {32'hc28a109c, 32'hc0e8103c} /* (6, 23, 10) {real, imag} */,
  {32'h41a6671f, 32'hc2ac1d82} /* (6, 23, 9) {real, imag} */,
  {32'hc2947597, 32'h424f47ac} /* (6, 23, 8) {real, imag} */,
  {32'hc1b0a85e, 32'h4275a488} /* (6, 23, 7) {real, imag} */,
  {32'hc1858e1b, 32'h42a6bbd3} /* (6, 23, 6) {real, imag} */,
  {32'hc2861237, 32'hc0552a80} /* (6, 23, 5) {real, imag} */,
  {32'h426166c0, 32'h422a60d8} /* (6, 23, 4) {real, imag} */,
  {32'h4229cce3, 32'h42eb0f83} /* (6, 23, 3) {real, imag} */,
  {32'hc4236a69, 32'hc2808a6a} /* (6, 23, 2) {real, imag} */,
  {32'h44afb9df, 32'h43cad4d7} /* (6, 23, 1) {real, imag} */,
  {32'h450ecaa4, 32'h00000000} /* (6, 23, 0) {real, imag} */,
  {32'h446f0367, 32'hc3ae6fd2} /* (6, 22, 31) {real, imag} */,
  {32'hc4331620, 32'h427a5af4} /* (6, 22, 30) {real, imag} */,
  {32'hc29be178, 32'hc3245b78} /* (6, 22, 29) {real, imag} */,
  {32'h4317eae2, 32'hc1da1ce8} /* (6, 22, 28) {real, imag} */,
  {32'hc281b8e6, 32'h430144be} /* (6, 22, 27) {real, imag} */,
  {32'h423f465c, 32'h419e4972} /* (6, 22, 26) {real, imag} */,
  {32'h42e99ec8, 32'hc24866d4} /* (6, 22, 25) {real, imag} */,
  {32'hc2a92df8, 32'h40909f00} /* (6, 22, 24) {real, imag} */,
  {32'hc2ec15fb, 32'hc166bb22} /* (6, 22, 23) {real, imag} */,
  {32'h42a5fceb, 32'hc2195e46} /* (6, 22, 22) {real, imag} */,
  {32'hbf8d3180, 32'h40b14948} /* (6, 22, 21) {real, imag} */,
  {32'h41b9e0f8, 32'hc16c9798} /* (6, 22, 20) {real, imag} */,
  {32'hc29b49be, 32'h427352cb} /* (6, 22, 19) {real, imag} */,
  {32'h4195f6e8, 32'h42388fe2} /* (6, 22, 18) {real, imag} */,
  {32'hc188c223, 32'hc194b424} /* (6, 22, 17) {real, imag} */,
  {32'hc203f83a, 32'h00000000} /* (6, 22, 16) {real, imag} */,
  {32'hc188c223, 32'h4194b424} /* (6, 22, 15) {real, imag} */,
  {32'h4195f6e8, 32'hc2388fe2} /* (6, 22, 14) {real, imag} */,
  {32'hc29b49be, 32'hc27352cb} /* (6, 22, 13) {real, imag} */,
  {32'h41b9e0f8, 32'h416c9798} /* (6, 22, 12) {real, imag} */,
  {32'hbf8d3180, 32'hc0b14948} /* (6, 22, 11) {real, imag} */,
  {32'h42a5fceb, 32'h42195e46} /* (6, 22, 10) {real, imag} */,
  {32'hc2ec15fb, 32'h4166bb22} /* (6, 22, 9) {real, imag} */,
  {32'hc2a92df8, 32'hc0909f00} /* (6, 22, 8) {real, imag} */,
  {32'h42e99ec8, 32'h424866d4} /* (6, 22, 7) {real, imag} */,
  {32'h423f465c, 32'hc19e4972} /* (6, 22, 6) {real, imag} */,
  {32'hc281b8e6, 32'hc30144be} /* (6, 22, 5) {real, imag} */,
  {32'h4317eae2, 32'h41da1ce8} /* (6, 22, 4) {real, imag} */,
  {32'hc29be178, 32'h43245b78} /* (6, 22, 3) {real, imag} */,
  {32'hc4331620, 32'hc27a5af4} /* (6, 22, 2) {real, imag} */,
  {32'h446f0367, 32'h43ae6fd2} /* (6, 22, 1) {real, imag} */,
  {32'h44e755a4, 32'h00000000} /* (6, 22, 0) {real, imag} */,
  {32'h43967708, 32'hc33b7084} /* (6, 21, 31) {real, imag} */,
  {32'hc3b67964, 32'hc310441f} /* (6, 21, 30) {real, imag} */,
  {32'hc3431ff5, 32'hc33963b1} /* (6, 21, 29) {real, imag} */,
  {32'hc171daf6, 32'h427944e3} /* (6, 21, 28) {real, imag} */,
  {32'h425b2c3e, 32'h42938c87} /* (6, 21, 27) {real, imag} */,
  {32'hc20b347c, 32'h42d0d68b} /* (6, 21, 26) {real, imag} */,
  {32'h428a7dc8, 32'h42bdc1d4} /* (6, 21, 25) {real, imag} */,
  {32'hc24cd535, 32'h41d0372b} /* (6, 21, 24) {real, imag} */,
  {32'h4227bcc6, 32'hbfb33d00} /* (6, 21, 23) {real, imag} */,
  {32'hc202514b, 32'hc286d99f} /* (6, 21, 22) {real, imag} */,
  {32'hc2596e28, 32'h4207d484} /* (6, 21, 21) {real, imag} */,
  {32'h41f3288a, 32'h42812890} /* (6, 21, 20) {real, imag} */,
  {32'h4209811e, 32'h428f08ed} /* (6, 21, 19) {real, imag} */,
  {32'hc1952762, 32'h418eab61} /* (6, 21, 18) {real, imag} */,
  {32'hc1c792ba, 32'hc3073cb8} /* (6, 21, 17) {real, imag} */,
  {32'h429d553a, 32'h00000000} /* (6, 21, 16) {real, imag} */,
  {32'hc1c792ba, 32'h43073cb8} /* (6, 21, 15) {real, imag} */,
  {32'hc1952762, 32'hc18eab61} /* (6, 21, 14) {real, imag} */,
  {32'h4209811e, 32'hc28f08ed} /* (6, 21, 13) {real, imag} */,
  {32'h41f3288a, 32'hc2812890} /* (6, 21, 12) {real, imag} */,
  {32'hc2596e28, 32'hc207d484} /* (6, 21, 11) {real, imag} */,
  {32'hc202514b, 32'h4286d99f} /* (6, 21, 10) {real, imag} */,
  {32'h4227bcc6, 32'h3fb33d00} /* (6, 21, 9) {real, imag} */,
  {32'hc24cd535, 32'hc1d0372b} /* (6, 21, 8) {real, imag} */,
  {32'h428a7dc8, 32'hc2bdc1d4} /* (6, 21, 7) {real, imag} */,
  {32'hc20b347c, 32'hc2d0d68b} /* (6, 21, 6) {real, imag} */,
  {32'h425b2c3e, 32'hc2938c87} /* (6, 21, 5) {real, imag} */,
  {32'hc171daf6, 32'hc27944e3} /* (6, 21, 4) {real, imag} */,
  {32'hc3431ff5, 32'h433963b1} /* (6, 21, 3) {real, imag} */,
  {32'hc3b67964, 32'h4310441f} /* (6, 21, 2) {real, imag} */,
  {32'h43967708, 32'h433b7084} /* (6, 21, 1) {real, imag} */,
  {32'h44a009c0, 32'h00000000} /* (6, 21, 0) {real, imag} */,
  {32'hc4430f92, 32'hc308aaf8} /* (6, 20, 31) {real, imag} */,
  {32'h43b9985c, 32'hc3386c8d} /* (6, 20, 30) {real, imag} */,
  {32'hc3323e9c, 32'hc315ee62} /* (6, 20, 29) {real, imag} */,
  {32'hc30bc4da, 32'hc2374b98} /* (6, 20, 28) {real, imag} */,
  {32'h42dedf7b, 32'hbfdd2ca0} /* (6, 20, 27) {real, imag} */,
  {32'hc186b3fe, 32'h421c4327} /* (6, 20, 26) {real, imag} */,
  {32'h41eacfa2, 32'h40a1e330} /* (6, 20, 25) {real, imag} */,
  {32'h41f75bcc, 32'hc07be8c8} /* (6, 20, 24) {real, imag} */,
  {32'hc26af5bf, 32'h42077cdd} /* (6, 20, 23) {real, imag} */,
  {32'hc2c40b66, 32'hc1a6d29c} /* (6, 20, 22) {real, imag} */,
  {32'h425817c0, 32'hc251c0ea} /* (6, 20, 21) {real, imag} */,
  {32'h422e0f3c, 32'hc00a0c20} /* (6, 20, 20) {real, imag} */,
  {32'hc19a01b4, 32'hc22f39b4} /* (6, 20, 19) {real, imag} */,
  {32'h4121a3f2, 32'hc179ebbc} /* (6, 20, 18) {real, imag} */,
  {32'h4268a809, 32'h42804a90} /* (6, 20, 17) {real, imag} */,
  {32'h42bc1498, 32'h00000000} /* (6, 20, 16) {real, imag} */,
  {32'h4268a809, 32'hc2804a90} /* (6, 20, 15) {real, imag} */,
  {32'h4121a3f2, 32'h4179ebbc} /* (6, 20, 14) {real, imag} */,
  {32'hc19a01b4, 32'h422f39b4} /* (6, 20, 13) {real, imag} */,
  {32'h422e0f3c, 32'h400a0c20} /* (6, 20, 12) {real, imag} */,
  {32'h425817c0, 32'h4251c0ea} /* (6, 20, 11) {real, imag} */,
  {32'hc2c40b66, 32'h41a6d29c} /* (6, 20, 10) {real, imag} */,
  {32'hc26af5bf, 32'hc2077cdd} /* (6, 20, 9) {real, imag} */,
  {32'h41f75bcc, 32'h407be8c8} /* (6, 20, 8) {real, imag} */,
  {32'h41eacfa2, 32'hc0a1e330} /* (6, 20, 7) {real, imag} */,
  {32'hc186b3fe, 32'hc21c4327} /* (6, 20, 6) {real, imag} */,
  {32'h42dedf7b, 32'h3fdd2ca0} /* (6, 20, 5) {real, imag} */,
  {32'hc30bc4da, 32'h42374b98} /* (6, 20, 4) {real, imag} */,
  {32'hc3323e9c, 32'h4315ee62} /* (6, 20, 3) {real, imag} */,
  {32'h43b9985c, 32'h43386c8d} /* (6, 20, 2) {real, imag} */,
  {32'hc4430f92, 32'h4308aaf8} /* (6, 20, 1) {real, imag} */,
  {32'h434b5c80, 32'h00000000} /* (6, 20, 0) {real, imag} */,
  {32'hc4b0c8e3, 32'h4353e210} /* (6, 19, 31) {real, imag} */,
  {32'h441dffa8, 32'hc2c13162} /* (6, 19, 30) {real, imag} */,
  {32'hc356c294, 32'hc39accd6} /* (6, 19, 29) {real, imag} */,
  {32'hc30185d8, 32'hc215b02b} /* (6, 19, 28) {real, imag} */,
  {32'h4302a388, 32'h40f87104} /* (6, 19, 27) {real, imag} */,
  {32'hc232f9ba, 32'h41c2cf7f} /* (6, 19, 26) {real, imag} */,
  {32'hc1709cdc, 32'hc2c72606} /* (6, 19, 25) {real, imag} */,
  {32'h41ec3e48, 32'hc19daaa5} /* (6, 19, 24) {real, imag} */,
  {32'hc28b4cba, 32'hc28bc5b8} /* (6, 19, 23) {real, imag} */,
  {32'h40f28ab8, 32'hc29677f5} /* (6, 19, 22) {real, imag} */,
  {32'h42e2bb12, 32'h419edd04} /* (6, 19, 21) {real, imag} */,
  {32'hc297289f, 32'h423c8846} /* (6, 19, 20) {real, imag} */,
  {32'hc15c8512, 32'hc1dcf4b8} /* (6, 19, 19) {real, imag} */,
  {32'h413ba174, 32'h41b91e00} /* (6, 19, 18) {real, imag} */,
  {32'h41a0c2a0, 32'hc0cdc088} /* (6, 19, 17) {real, imag} */,
  {32'h42031ea8, 32'h00000000} /* (6, 19, 16) {real, imag} */,
  {32'h41a0c2a0, 32'h40cdc088} /* (6, 19, 15) {real, imag} */,
  {32'h413ba174, 32'hc1b91e00} /* (6, 19, 14) {real, imag} */,
  {32'hc15c8512, 32'h41dcf4b8} /* (6, 19, 13) {real, imag} */,
  {32'hc297289f, 32'hc23c8846} /* (6, 19, 12) {real, imag} */,
  {32'h42e2bb12, 32'hc19edd04} /* (6, 19, 11) {real, imag} */,
  {32'h40f28ab8, 32'h429677f5} /* (6, 19, 10) {real, imag} */,
  {32'hc28b4cba, 32'h428bc5b8} /* (6, 19, 9) {real, imag} */,
  {32'h41ec3e48, 32'h419daaa5} /* (6, 19, 8) {real, imag} */,
  {32'hc1709cdc, 32'h42c72606} /* (6, 19, 7) {real, imag} */,
  {32'hc232f9ba, 32'hc1c2cf7f} /* (6, 19, 6) {real, imag} */,
  {32'h4302a388, 32'hc0f87104} /* (6, 19, 5) {real, imag} */,
  {32'hc30185d8, 32'h4215b02b} /* (6, 19, 4) {real, imag} */,
  {32'hc356c294, 32'h439accd6} /* (6, 19, 3) {real, imag} */,
  {32'h441dffa8, 32'h42c13162} /* (6, 19, 2) {real, imag} */,
  {32'hc4b0c8e3, 32'hc353e210} /* (6, 19, 1) {real, imag} */,
  {32'hc3d1a462, 32'h00000000} /* (6, 19, 0) {real, imag} */,
  {32'hc4e88566, 32'h4328dad7} /* (6, 18, 31) {real, imag} */,
  {32'h4446c93c, 32'hc19f0ef0} /* (6, 18, 30) {real, imag} */,
  {32'hc315fa3b, 32'hc331ab46} /* (6, 18, 29) {real, imag} */,
  {32'hc32e777b, 32'hc25f031a} /* (6, 18, 28) {real, imag} */,
  {32'h43215f31, 32'h41642d8c} /* (6, 18, 27) {real, imag} */,
  {32'h4295032a, 32'h4193dc97} /* (6, 18, 26) {real, imag} */,
  {32'h41844402, 32'h41f88235} /* (6, 18, 25) {real, imag} */,
  {32'hc2bd96d6, 32'h424c2222} /* (6, 18, 24) {real, imag} */,
  {32'hc215966d, 32'h411ecdd9} /* (6, 18, 23) {real, imag} */,
  {32'h42dd1f00, 32'h41314a54} /* (6, 18, 22) {real, imag} */,
  {32'hc21ae48d, 32'hc2a331a6} /* (6, 18, 21) {real, imag} */,
  {32'hc2a67722, 32'h41788cc4} /* (6, 18, 20) {real, imag} */,
  {32'h4227da53, 32'h41cc4f72} /* (6, 18, 19) {real, imag} */,
  {32'h42465e25, 32'hc1494614} /* (6, 18, 18) {real, imag} */,
  {32'h413383d6, 32'h4181d486} /* (6, 18, 17) {real, imag} */,
  {32'hc28b31d0, 32'h00000000} /* (6, 18, 16) {real, imag} */,
  {32'h413383d6, 32'hc181d486} /* (6, 18, 15) {real, imag} */,
  {32'h42465e25, 32'h41494614} /* (6, 18, 14) {real, imag} */,
  {32'h4227da53, 32'hc1cc4f72} /* (6, 18, 13) {real, imag} */,
  {32'hc2a67722, 32'hc1788cc4} /* (6, 18, 12) {real, imag} */,
  {32'hc21ae48d, 32'h42a331a6} /* (6, 18, 11) {real, imag} */,
  {32'h42dd1f00, 32'hc1314a54} /* (6, 18, 10) {real, imag} */,
  {32'hc215966d, 32'hc11ecdd9} /* (6, 18, 9) {real, imag} */,
  {32'hc2bd96d6, 32'hc24c2222} /* (6, 18, 8) {real, imag} */,
  {32'h41844402, 32'hc1f88235} /* (6, 18, 7) {real, imag} */,
  {32'h4295032a, 32'hc193dc97} /* (6, 18, 6) {real, imag} */,
  {32'h43215f31, 32'hc1642d8c} /* (6, 18, 5) {real, imag} */,
  {32'hc32e777b, 32'h425f031a} /* (6, 18, 4) {real, imag} */,
  {32'hc315fa3b, 32'h4331ab46} /* (6, 18, 3) {real, imag} */,
  {32'h4446c93c, 32'h419f0ef0} /* (6, 18, 2) {real, imag} */,
  {32'hc4e88566, 32'hc328dad7} /* (6, 18, 1) {real, imag} */,
  {32'hc43eafb1, 32'h00000000} /* (6, 18, 0) {real, imag} */,
  {32'hc503cdbf, 32'h430ad0bb} /* (6, 17, 31) {real, imag} */,
  {32'h44614028, 32'hc2ada668} /* (6, 17, 30) {real, imag} */,
  {32'hc2856265, 32'hc1ff83d8} /* (6, 17, 29) {real, imag} */,
  {32'hc2ea8e91, 32'hc23e9df4} /* (6, 17, 28) {real, imag} */,
  {32'h42d17cd5, 32'h42948515} /* (6, 17, 27) {real, imag} */,
  {32'h40a2fb48, 32'h42bcf1c6} /* (6, 17, 26) {real, imag} */,
  {32'h41229a86, 32'hc2cb5faa} /* (6, 17, 25) {real, imag} */,
  {32'h42e0791b, 32'hc2470049} /* (6, 17, 24) {real, imag} */,
  {32'hc26536d3, 32'h425b37ec} /* (6, 17, 23) {real, imag} */,
  {32'hc279c531, 32'h4262a2ce} /* (6, 17, 22) {real, imag} */,
  {32'h421a3b4a, 32'hc2a66a24} /* (6, 17, 21) {real, imag} */,
  {32'hc12475e4, 32'hc23ccd72} /* (6, 17, 20) {real, imag} */,
  {32'h4262ff0c, 32'h41886b07} /* (6, 17, 19) {real, imag} */,
  {32'hc25c6b0a, 32'h42254f1e} /* (6, 17, 18) {real, imag} */,
  {32'hc042e9e4, 32'hc234bc62} /* (6, 17, 17) {real, imag} */,
  {32'h420f8eab, 32'h00000000} /* (6, 17, 16) {real, imag} */,
  {32'hc042e9e4, 32'h4234bc62} /* (6, 17, 15) {real, imag} */,
  {32'hc25c6b0a, 32'hc2254f1e} /* (6, 17, 14) {real, imag} */,
  {32'h4262ff0c, 32'hc1886b07} /* (6, 17, 13) {real, imag} */,
  {32'hc12475e4, 32'h423ccd72} /* (6, 17, 12) {real, imag} */,
  {32'h421a3b4a, 32'h42a66a24} /* (6, 17, 11) {real, imag} */,
  {32'hc279c531, 32'hc262a2ce} /* (6, 17, 10) {real, imag} */,
  {32'hc26536d3, 32'hc25b37ec} /* (6, 17, 9) {real, imag} */,
  {32'h42e0791b, 32'h42470049} /* (6, 17, 8) {real, imag} */,
  {32'h41229a86, 32'h42cb5faa} /* (6, 17, 7) {real, imag} */,
  {32'h40a2fb48, 32'hc2bcf1c6} /* (6, 17, 6) {real, imag} */,
  {32'h42d17cd5, 32'hc2948515} /* (6, 17, 5) {real, imag} */,
  {32'hc2ea8e91, 32'h423e9df4} /* (6, 17, 4) {real, imag} */,
  {32'hc2856265, 32'h41ff83d8} /* (6, 17, 3) {real, imag} */,
  {32'h44614028, 32'h42ada668} /* (6, 17, 2) {real, imag} */,
  {32'hc503cdbf, 32'hc30ad0bb} /* (6, 17, 1) {real, imag} */,
  {32'hc490a38a, 32'h00000000} /* (6, 17, 0) {real, imag} */,
  {32'hc510a1d4, 32'h42300420} /* (6, 16, 31) {real, imag} */,
  {32'h444892b4, 32'hc34e9d43} /* (6, 16, 30) {real, imag} */,
  {32'hc2d7b351, 32'hc2226afe} /* (6, 16, 29) {real, imag} */,
  {32'hc29ea0b0, 32'hc2f2ae3e} /* (6, 16, 28) {real, imag} */,
  {32'h42ba71c6, 32'hc28af93a} /* (6, 16, 27) {real, imag} */,
  {32'h41d35f4a, 32'hc30e6d4e} /* (6, 16, 26) {real, imag} */,
  {32'h426b3f88, 32'h423f18b0} /* (6, 16, 25) {real, imag} */,
  {32'h42522916, 32'hc2d1b7ec} /* (6, 16, 24) {real, imag} */,
  {32'hc277d978, 32'hc29aaa48} /* (6, 16, 23) {real, imag} */,
  {32'h41337114, 32'hc302d09e} /* (6, 16, 22) {real, imag} */,
  {32'h4294c0f0, 32'hc252af6e} /* (6, 16, 21) {real, imag} */,
  {32'hc2295c10, 32'hc23b716e} /* (6, 16, 20) {real, imag} */,
  {32'h4184664c, 32'h42adadb4} /* (6, 16, 19) {real, imag} */,
  {32'h4115e430, 32'hbea81b00} /* (6, 16, 18) {real, imag} */,
  {32'h4259dc64, 32'hc2298518} /* (6, 16, 17) {real, imag} */,
  {32'h41dfd182, 32'h00000000} /* (6, 16, 16) {real, imag} */,
  {32'h4259dc64, 32'h42298518} /* (6, 16, 15) {real, imag} */,
  {32'h4115e430, 32'h3ea81b00} /* (6, 16, 14) {real, imag} */,
  {32'h4184664c, 32'hc2adadb4} /* (6, 16, 13) {real, imag} */,
  {32'hc2295c10, 32'h423b716e} /* (6, 16, 12) {real, imag} */,
  {32'h4294c0f0, 32'h4252af6e} /* (6, 16, 11) {real, imag} */,
  {32'h41337114, 32'h4302d09e} /* (6, 16, 10) {real, imag} */,
  {32'hc277d978, 32'h429aaa48} /* (6, 16, 9) {real, imag} */,
  {32'h42522916, 32'h42d1b7ec} /* (6, 16, 8) {real, imag} */,
  {32'h426b3f88, 32'hc23f18b0} /* (6, 16, 7) {real, imag} */,
  {32'h41d35f4a, 32'h430e6d4e} /* (6, 16, 6) {real, imag} */,
  {32'h42ba71c6, 32'h428af93a} /* (6, 16, 5) {real, imag} */,
  {32'hc29ea0b0, 32'h42f2ae3e} /* (6, 16, 4) {real, imag} */,
  {32'hc2d7b351, 32'h42226afe} /* (6, 16, 3) {real, imag} */,
  {32'h444892b4, 32'h434e9d43} /* (6, 16, 2) {real, imag} */,
  {32'hc510a1d4, 32'hc2300420} /* (6, 16, 1) {real, imag} */,
  {32'hc4cf5ba8, 32'h00000000} /* (6, 16, 0) {real, imag} */,
  {32'hc50ce4c5, 32'hc10b8d30} /* (6, 15, 31) {real, imag} */,
  {32'h444353c4, 32'hc30955b8} /* (6, 15, 30) {real, imag} */,
  {32'hc1d1dd54, 32'hc326253f} /* (6, 15, 29) {real, imag} */,
  {32'hc3175b5d, 32'hc3503e71} /* (6, 15, 28) {real, imag} */,
  {32'h429e390f, 32'hc2f664c5} /* (6, 15, 27) {real, imag} */,
  {32'h42f97580, 32'hc355e289} /* (6, 15, 26) {real, imag} */,
  {32'h42899bc9, 32'h42533087} /* (6, 15, 25) {real, imag} */,
  {32'h428af1bf, 32'hc20ebccf} /* (6, 15, 24) {real, imag} */,
  {32'hc284f549, 32'h41988f00} /* (6, 15, 23) {real, imag} */,
  {32'h42b6333c, 32'h41c8ae40} /* (6, 15, 22) {real, imag} */,
  {32'hc09ece2c, 32'hc27170c9} /* (6, 15, 21) {real, imag} */,
  {32'h4246816f, 32'hc2ad3c2d} /* (6, 15, 20) {real, imag} */,
  {32'hc2679e70, 32'hc1f33cf5} /* (6, 15, 19) {real, imag} */,
  {32'hc21ee12a, 32'h40eb7394} /* (6, 15, 18) {real, imag} */,
  {32'hc1b553ac, 32'h4254ccb2} /* (6, 15, 17) {real, imag} */,
  {32'h42a49848, 32'h00000000} /* (6, 15, 16) {real, imag} */,
  {32'hc1b553ac, 32'hc254ccb2} /* (6, 15, 15) {real, imag} */,
  {32'hc21ee12a, 32'hc0eb7394} /* (6, 15, 14) {real, imag} */,
  {32'hc2679e70, 32'h41f33cf5} /* (6, 15, 13) {real, imag} */,
  {32'h4246816f, 32'h42ad3c2d} /* (6, 15, 12) {real, imag} */,
  {32'hc09ece2c, 32'h427170c9} /* (6, 15, 11) {real, imag} */,
  {32'h42b6333c, 32'hc1c8ae40} /* (6, 15, 10) {real, imag} */,
  {32'hc284f549, 32'hc1988f00} /* (6, 15, 9) {real, imag} */,
  {32'h428af1bf, 32'h420ebccf} /* (6, 15, 8) {real, imag} */,
  {32'h42899bc9, 32'hc2533087} /* (6, 15, 7) {real, imag} */,
  {32'h42f97580, 32'h4355e289} /* (6, 15, 6) {real, imag} */,
  {32'h429e390f, 32'h42f664c5} /* (6, 15, 5) {real, imag} */,
  {32'hc3175b5d, 32'h43503e71} /* (6, 15, 4) {real, imag} */,
  {32'hc1d1dd54, 32'h4326253f} /* (6, 15, 3) {real, imag} */,
  {32'h444353c4, 32'h430955b8} /* (6, 15, 2) {real, imag} */,
  {32'hc50ce4c5, 32'h410b8d30} /* (6, 15, 1) {real, imag} */,
  {32'hc4de820a, 32'h00000000} /* (6, 15, 0) {real, imag} */,
  {32'hc4f08f4e, 32'h42507204} /* (6, 14, 31) {real, imag} */,
  {32'h44688a4a, 32'hc2f4db34} /* (6, 14, 30) {real, imag} */,
  {32'h422c0a00, 32'hc2821ed4} /* (6, 14, 29) {real, imag} */,
  {32'hc3246699, 32'hc328b4c8} /* (6, 14, 28) {real, imag} */,
  {32'h432a79cb, 32'h4273208f} /* (6, 14, 27) {real, imag} */,
  {32'h425e6644, 32'hc29bbb0a} /* (6, 14, 26) {real, imag} */,
  {32'hc1d95bf6, 32'hc289642b} /* (6, 14, 25) {real, imag} */,
  {32'h43393d59, 32'hc00120d8} /* (6, 14, 24) {real, imag} */,
  {32'h41f1abaa, 32'h4193cc44} /* (6, 14, 23) {real, imag} */,
  {32'hc2c3bbcc, 32'h42a9eb26} /* (6, 14, 22) {real, imag} */,
  {32'h42099933, 32'hc1f0e01a} /* (6, 14, 21) {real, imag} */,
  {32'h42d0accc, 32'h42bf06e4} /* (6, 14, 20) {real, imag} */,
  {32'hc217d167, 32'h41911622} /* (6, 14, 19) {real, imag} */,
  {32'hc102c754, 32'hc2a4b28e} /* (6, 14, 18) {real, imag} */,
  {32'hc27c9aa6, 32'h42936a40} /* (6, 14, 17) {real, imag} */,
  {32'hc0518250, 32'h00000000} /* (6, 14, 16) {real, imag} */,
  {32'hc27c9aa6, 32'hc2936a40} /* (6, 14, 15) {real, imag} */,
  {32'hc102c754, 32'h42a4b28e} /* (6, 14, 14) {real, imag} */,
  {32'hc217d167, 32'hc1911622} /* (6, 14, 13) {real, imag} */,
  {32'h42d0accc, 32'hc2bf06e4} /* (6, 14, 12) {real, imag} */,
  {32'h42099933, 32'h41f0e01a} /* (6, 14, 11) {real, imag} */,
  {32'hc2c3bbcc, 32'hc2a9eb26} /* (6, 14, 10) {real, imag} */,
  {32'h41f1abaa, 32'hc193cc44} /* (6, 14, 9) {real, imag} */,
  {32'h43393d59, 32'h400120d8} /* (6, 14, 8) {real, imag} */,
  {32'hc1d95bf6, 32'h4289642b} /* (6, 14, 7) {real, imag} */,
  {32'h425e6644, 32'h429bbb0a} /* (6, 14, 6) {real, imag} */,
  {32'h432a79cb, 32'hc273208f} /* (6, 14, 5) {real, imag} */,
  {32'hc3246699, 32'h4328b4c8} /* (6, 14, 4) {real, imag} */,
  {32'h422c0a00, 32'h42821ed4} /* (6, 14, 3) {real, imag} */,
  {32'h44688a4a, 32'h42f4db34} /* (6, 14, 2) {real, imag} */,
  {32'hc4f08f4e, 32'hc2507204} /* (6, 14, 1) {real, imag} */,
  {32'hc4e249ce, 32'h00000000} /* (6, 14, 0) {real, imag} */,
  {32'hc4c8675b, 32'hc226efc0} /* (6, 13, 31) {real, imag} */,
  {32'h446f3c68, 32'hc30a5315} /* (6, 13, 30) {real, imag} */,
  {32'h429856bc, 32'h420e127c} /* (6, 13, 29) {real, imag} */,
  {32'hc31521c8, 32'hc2a691c4} /* (6, 13, 28) {real, imag} */,
  {32'h437711e0, 32'h41261e4a} /* (6, 13, 27) {real, imag} */,
  {32'h42fd9317, 32'h4275c632} /* (6, 13, 26) {real, imag} */,
  {32'hc20d53f8, 32'hc27bda43} /* (6, 13, 25) {real, imag} */,
  {32'h430bfe43, 32'h415d6f2a} /* (6, 13, 24) {real, imag} */,
  {32'hc22a9a0b, 32'h433f31ee} /* (6, 13, 23) {real, imag} */,
  {32'hc2b55da4, 32'h42ab16c1} /* (6, 13, 22) {real, imag} */,
  {32'h41ca123a, 32'hc3545cf4} /* (6, 13, 21) {real, imag} */,
  {32'h41afb1bc, 32'hc2c2cda5} /* (6, 13, 20) {real, imag} */,
  {32'h41c499b5, 32'h43398ed2} /* (6, 13, 19) {real, imag} */,
  {32'hc26cd3bf, 32'hc2e4cf30} /* (6, 13, 18) {real, imag} */,
  {32'h4283537c, 32'hc104c20a} /* (6, 13, 17) {real, imag} */,
  {32'h4174be8e, 32'h00000000} /* (6, 13, 16) {real, imag} */,
  {32'h4283537c, 32'h4104c20a} /* (6, 13, 15) {real, imag} */,
  {32'hc26cd3bf, 32'h42e4cf30} /* (6, 13, 14) {real, imag} */,
  {32'h41c499b5, 32'hc3398ed2} /* (6, 13, 13) {real, imag} */,
  {32'h41afb1bc, 32'h42c2cda5} /* (6, 13, 12) {real, imag} */,
  {32'h41ca123a, 32'h43545cf4} /* (6, 13, 11) {real, imag} */,
  {32'hc2b55da4, 32'hc2ab16c1} /* (6, 13, 10) {real, imag} */,
  {32'hc22a9a0b, 32'hc33f31ee} /* (6, 13, 9) {real, imag} */,
  {32'h430bfe43, 32'hc15d6f2a} /* (6, 13, 8) {real, imag} */,
  {32'hc20d53f8, 32'h427bda43} /* (6, 13, 7) {real, imag} */,
  {32'h42fd9317, 32'hc275c632} /* (6, 13, 6) {real, imag} */,
  {32'h437711e0, 32'hc1261e4a} /* (6, 13, 5) {real, imag} */,
  {32'hc31521c8, 32'h42a691c4} /* (6, 13, 4) {real, imag} */,
  {32'h429856bc, 32'hc20e127c} /* (6, 13, 3) {real, imag} */,
  {32'h446f3c68, 32'h430a5315} /* (6, 13, 2) {real, imag} */,
  {32'hc4c8675b, 32'h4226efc0} /* (6, 13, 1) {real, imag} */,
  {32'hc4cdbb32, 32'h00000000} /* (6, 13, 0) {real, imag} */,
  {32'hc4968af1, 32'hc14f7500} /* (6, 12, 31) {real, imag} */,
  {32'h443475ac, 32'hc349c0fb} /* (6, 12, 30) {real, imag} */,
  {32'h4306abee, 32'h4274799c} /* (6, 12, 29) {real, imag} */,
  {32'hc345d97a, 32'hc23df7a4} /* (6, 12, 28) {real, imag} */,
  {32'h42cb6f61, 32'hc20627f9} /* (6, 12, 27) {real, imag} */,
  {32'h4265e1b9, 32'h43040f20} /* (6, 12, 26) {real, imag} */,
  {32'hc197494a, 32'hc2aba2b3} /* (6, 12, 25) {real, imag} */,
  {32'h42ef2b0b, 32'h41517aae} /* (6, 12, 24) {real, imag} */,
  {32'hc23176d3, 32'hc06f8850} /* (6, 12, 23) {real, imag} */,
  {32'h4302c4bc, 32'hc2528eaa} /* (6, 12, 22) {real, imag} */,
  {32'hc0534d58, 32'h4121cb5a} /* (6, 12, 21) {real, imag} */,
  {32'hc2f9d8d6, 32'h426f79fb} /* (6, 12, 20) {real, imag} */,
  {32'h42ea3873, 32'hc2dc1df2} /* (6, 12, 19) {real, imag} */,
  {32'h3fec5570, 32'h4207953f} /* (6, 12, 18) {real, imag} */,
  {32'hc26432eb, 32'h4205383c} /* (6, 12, 17) {real, imag} */,
  {32'h4181bf6a, 32'h00000000} /* (6, 12, 16) {real, imag} */,
  {32'hc26432eb, 32'hc205383c} /* (6, 12, 15) {real, imag} */,
  {32'h3fec5570, 32'hc207953f} /* (6, 12, 14) {real, imag} */,
  {32'h42ea3873, 32'h42dc1df2} /* (6, 12, 13) {real, imag} */,
  {32'hc2f9d8d6, 32'hc26f79fb} /* (6, 12, 12) {real, imag} */,
  {32'hc0534d58, 32'hc121cb5a} /* (6, 12, 11) {real, imag} */,
  {32'h4302c4bc, 32'h42528eaa} /* (6, 12, 10) {real, imag} */,
  {32'hc23176d3, 32'h406f8850} /* (6, 12, 9) {real, imag} */,
  {32'h42ef2b0b, 32'hc1517aae} /* (6, 12, 8) {real, imag} */,
  {32'hc197494a, 32'h42aba2b3} /* (6, 12, 7) {real, imag} */,
  {32'h4265e1b9, 32'hc3040f20} /* (6, 12, 6) {real, imag} */,
  {32'h42cb6f61, 32'h420627f9} /* (6, 12, 5) {real, imag} */,
  {32'hc345d97a, 32'h423df7a4} /* (6, 12, 4) {real, imag} */,
  {32'h4306abee, 32'hc274799c} /* (6, 12, 3) {real, imag} */,
  {32'h443475ac, 32'h4349c0fb} /* (6, 12, 2) {real, imag} */,
  {32'hc4968af1, 32'h414f7500} /* (6, 12, 1) {real, imag} */,
  {32'hc47a979c, 32'h00000000} /* (6, 12, 0) {real, imag} */,
  {32'hc42142a8, 32'hc3856d56} /* (6, 11, 31) {real, imag} */,
  {32'h43fe04e8, 32'hc2f136e6} /* (6, 11, 30) {real, imag} */,
  {32'h4352fe07, 32'h4294812a} /* (6, 11, 29) {real, imag} */,
  {32'hc075f668, 32'hc2c18172} /* (6, 11, 28) {real, imag} */,
  {32'h428cfd52, 32'hc28f642b} /* (6, 11, 27) {real, imag} */,
  {32'hc13068c9, 32'h4249444e} /* (6, 11, 26) {real, imag} */,
  {32'hc238edff, 32'hc2bb209e} /* (6, 11, 25) {real, imag} */,
  {32'h3f143080, 32'hc2b240ad} /* (6, 11, 24) {real, imag} */,
  {32'h41fa6ebc, 32'hc2d4efb7} /* (6, 11, 23) {real, imag} */,
  {32'h41e96ca6, 32'h4295bae9} /* (6, 11, 22) {real, imag} */,
  {32'h401fb980, 32'hc1fa1210} /* (6, 11, 21) {real, imag} */,
  {32'h41d9839a, 32'h4269e704} /* (6, 11, 20) {real, imag} */,
  {32'h419f0af5, 32'h425dd9fa} /* (6, 11, 19) {real, imag} */,
  {32'h413a9dcc, 32'h423e08de} /* (6, 11, 18) {real, imag} */,
  {32'hc166c203, 32'h42245f7a} /* (6, 11, 17) {real, imag} */,
  {32'h41dfeaa7, 32'h00000000} /* (6, 11, 16) {real, imag} */,
  {32'hc166c203, 32'hc2245f7a} /* (6, 11, 15) {real, imag} */,
  {32'h413a9dcc, 32'hc23e08de} /* (6, 11, 14) {real, imag} */,
  {32'h419f0af5, 32'hc25dd9fa} /* (6, 11, 13) {real, imag} */,
  {32'h41d9839a, 32'hc269e704} /* (6, 11, 12) {real, imag} */,
  {32'h401fb980, 32'h41fa1210} /* (6, 11, 11) {real, imag} */,
  {32'h41e96ca6, 32'hc295bae9} /* (6, 11, 10) {real, imag} */,
  {32'h41fa6ebc, 32'h42d4efb7} /* (6, 11, 9) {real, imag} */,
  {32'h3f143080, 32'h42b240ad} /* (6, 11, 8) {real, imag} */,
  {32'hc238edff, 32'h42bb209e} /* (6, 11, 7) {real, imag} */,
  {32'hc13068c9, 32'hc249444e} /* (6, 11, 6) {real, imag} */,
  {32'h428cfd52, 32'h428f642b} /* (6, 11, 5) {real, imag} */,
  {32'hc075f668, 32'h42c18172} /* (6, 11, 4) {real, imag} */,
  {32'h4352fe07, 32'hc294812a} /* (6, 11, 3) {real, imag} */,
  {32'h43fe04e8, 32'h42f136e6} /* (6, 11, 2) {real, imag} */,
  {32'hc42142a8, 32'h43856d56} /* (6, 11, 1) {real, imag} */,
  {32'hc4039db1, 32'h00000000} /* (6, 11, 0) {real, imag} */,
  {32'h43ecafc6, 32'hc404e303} /* (6, 10, 31) {real, imag} */,
  {32'hc2da882c, 32'h422ee31c} /* (6, 10, 30) {real, imag} */,
  {32'h42892cb4, 32'h427d150a} /* (6, 10, 29) {real, imag} */,
  {32'h42a1f2fd, 32'hc3530961} /* (6, 10, 28) {real, imag} */,
  {32'hc1bbc521, 32'h429f5f95} /* (6, 10, 27) {real, imag} */,
  {32'h41ea6280, 32'h425cfc03} /* (6, 10, 26) {real, imag} */,
  {32'h42af1b68, 32'h41699bc2} /* (6, 10, 25) {real, imag} */,
  {32'h4229edb7, 32'h4224974e} /* (6, 10, 24) {real, imag} */,
  {32'h42d7dcff, 32'hc220a17e} /* (6, 10, 23) {real, imag} */,
  {32'hc2202838, 32'hc23a26aa} /* (6, 10, 22) {real, imag} */,
  {32'hc1611298, 32'h42d2a1f0} /* (6, 10, 21) {real, imag} */,
  {32'hc27491bc, 32'h41932658} /* (6, 10, 20) {real, imag} */,
  {32'hc18c005b, 32'h420f45d3} /* (6, 10, 19) {real, imag} */,
  {32'h427cea6e, 32'hc20d1aca} /* (6, 10, 18) {real, imag} */,
  {32'hc18d68e7, 32'h4266de1a} /* (6, 10, 17) {real, imag} */,
  {32'h40428718, 32'h00000000} /* (6, 10, 16) {real, imag} */,
  {32'hc18d68e7, 32'hc266de1a} /* (6, 10, 15) {real, imag} */,
  {32'h427cea6e, 32'h420d1aca} /* (6, 10, 14) {real, imag} */,
  {32'hc18c005b, 32'hc20f45d3} /* (6, 10, 13) {real, imag} */,
  {32'hc27491bc, 32'hc1932658} /* (6, 10, 12) {real, imag} */,
  {32'hc1611298, 32'hc2d2a1f0} /* (6, 10, 11) {real, imag} */,
  {32'hc2202838, 32'h423a26aa} /* (6, 10, 10) {real, imag} */,
  {32'h42d7dcff, 32'h4220a17e} /* (6, 10, 9) {real, imag} */,
  {32'h4229edb7, 32'hc224974e} /* (6, 10, 8) {real, imag} */,
  {32'h42af1b68, 32'hc1699bc2} /* (6, 10, 7) {real, imag} */,
  {32'h41ea6280, 32'hc25cfc03} /* (6, 10, 6) {real, imag} */,
  {32'hc1bbc521, 32'hc29f5f95} /* (6, 10, 5) {real, imag} */,
  {32'h42a1f2fd, 32'h43530961} /* (6, 10, 4) {real, imag} */,
  {32'h42892cb4, 32'hc27d150a} /* (6, 10, 3) {real, imag} */,
  {32'hc2da882c, 32'hc22ee31c} /* (6, 10, 2) {real, imag} */,
  {32'h43ecafc6, 32'h4404e303} /* (6, 10, 1) {real, imag} */,
  {32'h442b821b, 32'h00000000} /* (6, 10, 0) {real, imag} */,
  {32'h449527e9, 32'hc437bd18} /* (6, 9, 31) {real, imag} */,
  {32'hc3e1d09e, 32'h4356fdd7} /* (6, 9, 30) {real, imag} */,
  {32'h42b389de, 32'h42887795} /* (6, 9, 29) {real, imag} */,
  {32'h42eb2a1e, 32'hc381aee9} /* (6, 9, 28) {real, imag} */,
  {32'hc2ae70ed, 32'h433ce4bf} /* (6, 9, 27) {real, imag} */,
  {32'hc2921251, 32'h42f53e09} /* (6, 9, 26) {real, imag} */,
  {32'h3e2b4340, 32'hc34100b6} /* (6, 9, 25) {real, imag} */,
  {32'hc312707e, 32'hc2d2ca78} /* (6, 9, 24) {real, imag} */,
  {32'hc1786496, 32'h42e1cece} /* (6, 9, 23) {real, imag} */,
  {32'hc2156adb, 32'hc21b1cce} /* (6, 9, 22) {real, imag} */,
  {32'hc2b2477e, 32'h433099b7} /* (6, 9, 21) {real, imag} */,
  {32'h41e810d3, 32'hc287e9fc} /* (6, 9, 20) {real, imag} */,
  {32'h4259e21c, 32'hc0bce324} /* (6, 9, 19) {real, imag} */,
  {32'h42d1532a, 32'h41d9d924} /* (6, 9, 18) {real, imag} */,
  {32'hc15bbc24, 32'hc29649e8} /* (6, 9, 17) {real, imag} */,
  {32'hc29a0d0e, 32'h00000000} /* (6, 9, 16) {real, imag} */,
  {32'hc15bbc24, 32'h429649e8} /* (6, 9, 15) {real, imag} */,
  {32'h42d1532a, 32'hc1d9d924} /* (6, 9, 14) {real, imag} */,
  {32'h4259e21c, 32'h40bce324} /* (6, 9, 13) {real, imag} */,
  {32'h41e810d3, 32'h4287e9fc} /* (6, 9, 12) {real, imag} */,
  {32'hc2b2477e, 32'hc33099b7} /* (6, 9, 11) {real, imag} */,
  {32'hc2156adb, 32'h421b1cce} /* (6, 9, 10) {real, imag} */,
  {32'hc1786496, 32'hc2e1cece} /* (6, 9, 9) {real, imag} */,
  {32'hc312707e, 32'h42d2ca78} /* (6, 9, 8) {real, imag} */,
  {32'h3e2b4340, 32'h434100b6} /* (6, 9, 7) {real, imag} */,
  {32'hc2921251, 32'hc2f53e09} /* (6, 9, 6) {real, imag} */,
  {32'hc2ae70ed, 32'hc33ce4bf} /* (6, 9, 5) {real, imag} */,
  {32'h42eb2a1e, 32'h4381aee9} /* (6, 9, 4) {real, imag} */,
  {32'h42b389de, 32'hc2887795} /* (6, 9, 3) {real, imag} */,
  {32'hc3e1d09e, 32'hc356fdd7} /* (6, 9, 2) {real, imag} */,
  {32'h449527e9, 32'h4437bd18} /* (6, 9, 1) {real, imag} */,
  {32'h44c6cd63, 32'h00000000} /* (6, 9, 0) {real, imag} */,
  {32'h44c105c7, 32'hc43d0352} /* (6, 8, 31) {real, imag} */,
  {32'hc3da60a2, 32'h43caf21a} /* (6, 8, 30) {real, imag} */,
  {32'h435776f1, 32'hc1bbe80c} /* (6, 8, 29) {real, imag} */,
  {32'h42bb21a4, 32'hc2eb378a} /* (6, 8, 28) {real, imag} */,
  {32'hc2f0757c, 32'h42a3eb70} /* (6, 8, 27) {real, imag} */,
  {32'hc2a3e665, 32'h42af30b7} /* (6, 8, 26) {real, imag} */,
  {32'hc2554abc, 32'hc2e7d9fc} /* (6, 8, 25) {real, imag} */,
  {32'hc2f6aa9b, 32'hc2c0fc9f} /* (6, 8, 24) {real, imag} */,
  {32'h42083394, 32'h4282430d} /* (6, 8, 23) {real, imag} */,
  {32'h41a93342, 32'h423c5360} /* (6, 8, 22) {real, imag} */,
  {32'h42898094, 32'h42de8655} /* (6, 8, 21) {real, imag} */,
  {32'h41e3a085, 32'h417ff398} /* (6, 8, 20) {real, imag} */,
  {32'h42923970, 32'h42255148} /* (6, 8, 19) {real, imag} */,
  {32'hc1bef1f9, 32'h4243ea45} /* (6, 8, 18) {real, imag} */,
  {32'h4206fb22, 32'hc1808e35} /* (6, 8, 17) {real, imag} */,
  {32'h4239fbad, 32'h00000000} /* (6, 8, 16) {real, imag} */,
  {32'h4206fb22, 32'h41808e35} /* (6, 8, 15) {real, imag} */,
  {32'hc1bef1f9, 32'hc243ea45} /* (6, 8, 14) {real, imag} */,
  {32'h42923970, 32'hc2255148} /* (6, 8, 13) {real, imag} */,
  {32'h41e3a085, 32'hc17ff398} /* (6, 8, 12) {real, imag} */,
  {32'h42898094, 32'hc2de8655} /* (6, 8, 11) {real, imag} */,
  {32'h41a93342, 32'hc23c5360} /* (6, 8, 10) {real, imag} */,
  {32'h42083394, 32'hc282430d} /* (6, 8, 9) {real, imag} */,
  {32'hc2f6aa9b, 32'h42c0fc9f} /* (6, 8, 8) {real, imag} */,
  {32'hc2554abc, 32'h42e7d9fc} /* (6, 8, 7) {real, imag} */,
  {32'hc2a3e665, 32'hc2af30b7} /* (6, 8, 6) {real, imag} */,
  {32'hc2f0757c, 32'hc2a3eb70} /* (6, 8, 5) {real, imag} */,
  {32'h42bb21a4, 32'h42eb378a} /* (6, 8, 4) {real, imag} */,
  {32'h435776f1, 32'h41bbe80c} /* (6, 8, 3) {real, imag} */,
  {32'hc3da60a2, 32'hc3caf21a} /* (6, 8, 2) {real, imag} */,
  {32'h44c105c7, 32'h443d0352} /* (6, 8, 1) {real, imag} */,
  {32'h44f67237, 32'h00000000} /* (6, 8, 0) {real, imag} */,
  {32'h44e54f2f, 32'hc4703c84} /* (6, 7, 31) {real, imag} */,
  {32'hc3fea696, 32'h441cd6e2} /* (6, 7, 30) {real, imag} */,
  {32'h437f176f, 32'hc1c21012} /* (6, 7, 29) {real, imag} */,
  {32'h42991d3b, 32'h40349330} /* (6, 7, 28) {real, imag} */,
  {32'hc32a16d9, 32'h40d767c0} /* (6, 7, 27) {real, imag} */,
  {32'h4171361e, 32'h3d38d800} /* (6, 7, 26) {real, imag} */,
  {32'h412ac34b, 32'hc2a865e8} /* (6, 7, 25) {real, imag} */,
  {32'hc2966855, 32'hc17f2b20} /* (6, 7, 24) {real, imag} */,
  {32'hc1ac54c3, 32'h4121c190} /* (6, 7, 23) {real, imag} */,
  {32'hc2bf9f5e, 32'hc2729fcd} /* (6, 7, 22) {real, imag} */,
  {32'h41bee6ec, 32'hc2814ed8} /* (6, 7, 21) {real, imag} */,
  {32'h41e6aff3, 32'hbf8e9460} /* (6, 7, 20) {real, imag} */,
  {32'hc225ea1a, 32'hc156ff82} /* (6, 7, 19) {real, imag} */,
  {32'hc1bc00a2, 32'h41d05e46} /* (6, 7, 18) {real, imag} */,
  {32'h4110c540, 32'hc124ef00} /* (6, 7, 17) {real, imag} */,
  {32'h428b8ef9, 32'h00000000} /* (6, 7, 16) {real, imag} */,
  {32'h4110c540, 32'h4124ef00} /* (6, 7, 15) {real, imag} */,
  {32'hc1bc00a2, 32'hc1d05e46} /* (6, 7, 14) {real, imag} */,
  {32'hc225ea1a, 32'h4156ff82} /* (6, 7, 13) {real, imag} */,
  {32'h41e6aff3, 32'h3f8e9460} /* (6, 7, 12) {real, imag} */,
  {32'h41bee6ec, 32'h42814ed8} /* (6, 7, 11) {real, imag} */,
  {32'hc2bf9f5e, 32'h42729fcd} /* (6, 7, 10) {real, imag} */,
  {32'hc1ac54c3, 32'hc121c190} /* (6, 7, 9) {real, imag} */,
  {32'hc2966855, 32'h417f2b20} /* (6, 7, 8) {real, imag} */,
  {32'h412ac34b, 32'h42a865e8} /* (6, 7, 7) {real, imag} */,
  {32'h4171361e, 32'hbd38d800} /* (6, 7, 6) {real, imag} */,
  {32'hc32a16d9, 32'hc0d767c0} /* (6, 7, 5) {real, imag} */,
  {32'h42991d3b, 32'hc0349330} /* (6, 7, 4) {real, imag} */,
  {32'h437f176f, 32'h41c21012} /* (6, 7, 3) {real, imag} */,
  {32'hc3fea696, 32'hc41cd6e2} /* (6, 7, 2) {real, imag} */,
  {32'h44e54f2f, 32'h44703c84} /* (6, 7, 1) {real, imag} */,
  {32'h45101a8c, 32'h00000000} /* (6, 7, 0) {real, imag} */,
  {32'h44fd7eb4, 32'hc471fe21} /* (6, 6, 31) {real, imag} */,
  {32'hc404cbee, 32'h4413635f} /* (6, 6, 30) {real, imag} */,
  {32'h4187cf68, 32'h3e40e800} /* (6, 6, 29) {real, imag} */,
  {32'h428c4ba1, 32'hc2e171dc} /* (6, 6, 28) {real, imag} */,
  {32'hc31010e7, 32'hc0f3d2d0} /* (6, 6, 27) {real, imag} */,
  {32'h429bf713, 32'hc1fea8a0} /* (6, 6, 26) {real, imag} */,
  {32'h42e6dbdd, 32'h4182f078} /* (6, 6, 25) {real, imag} */,
  {32'hc2cb7bf4, 32'h42dd2715} /* (6, 6, 24) {real, imag} */,
  {32'hc25ed971, 32'h41df948b} /* (6, 6, 23) {real, imag} */,
  {32'hc214b806, 32'h429b7b1d} /* (6, 6, 22) {real, imag} */,
  {32'hc2c9930c, 32'h422c1ebe} /* (6, 6, 21) {real, imag} */,
  {32'h430c35c6, 32'hc22ad735} /* (6, 6, 20) {real, imag} */,
  {32'h406dfad8, 32'hc250ef7f} /* (6, 6, 19) {real, imag} */,
  {32'hc1eb4646, 32'hc147a23e} /* (6, 6, 18) {real, imag} */,
  {32'h41afbc5d, 32'hc2052e74} /* (6, 6, 17) {real, imag} */,
  {32'hc0d5005e, 32'h00000000} /* (6, 6, 16) {real, imag} */,
  {32'h41afbc5d, 32'h42052e74} /* (6, 6, 15) {real, imag} */,
  {32'hc1eb4646, 32'h4147a23e} /* (6, 6, 14) {real, imag} */,
  {32'h406dfad8, 32'h4250ef7f} /* (6, 6, 13) {real, imag} */,
  {32'h430c35c6, 32'h422ad735} /* (6, 6, 12) {real, imag} */,
  {32'hc2c9930c, 32'hc22c1ebe} /* (6, 6, 11) {real, imag} */,
  {32'hc214b806, 32'hc29b7b1d} /* (6, 6, 10) {real, imag} */,
  {32'hc25ed971, 32'hc1df948b} /* (6, 6, 9) {real, imag} */,
  {32'hc2cb7bf4, 32'hc2dd2715} /* (6, 6, 8) {real, imag} */,
  {32'h42e6dbdd, 32'hc182f078} /* (6, 6, 7) {real, imag} */,
  {32'h429bf713, 32'h41fea8a0} /* (6, 6, 6) {real, imag} */,
  {32'hc31010e7, 32'h40f3d2d0} /* (6, 6, 5) {real, imag} */,
  {32'h428c4ba1, 32'h42e171dc} /* (6, 6, 4) {real, imag} */,
  {32'h4187cf68, 32'hbe40e800} /* (6, 6, 3) {real, imag} */,
  {32'hc404cbee, 32'hc413635f} /* (6, 6, 2) {real, imag} */,
  {32'h44fd7eb4, 32'h4471fe21} /* (6, 6, 1) {real, imag} */,
  {32'h4533946c, 32'h00000000} /* (6, 6, 0) {real, imag} */,
  {32'h44efa338, 32'hc4c32180} /* (6, 5, 31) {real, imag} */,
  {32'hc31cc9c4, 32'h4420e3ca} /* (6, 5, 30) {real, imag} */,
  {32'h41e28a5c, 32'h426a9ae3} /* (6, 5, 29) {real, imag} */,
  {32'h41cab508, 32'h4095f160} /* (6, 5, 28) {real, imag} */,
  {32'hc2ec9173, 32'hc2b9705b} /* (6, 5, 27) {real, imag} */,
  {32'h425e7127, 32'hc0bc862c} /* (6, 5, 26) {real, imag} */,
  {32'h42869de8, 32'hc29d56c4} /* (6, 5, 25) {real, imag} */,
  {32'hc09ddfb8, 32'hc17d5c52} /* (6, 5, 24) {real, imag} */,
  {32'hc2d084f6, 32'hc2f1d38e} /* (6, 5, 23) {real, imag} */,
  {32'h43131105, 32'hc22bd33b} /* (6, 5, 22) {real, imag} */,
  {32'hc2b7f392, 32'h42859a0b} /* (6, 5, 21) {real, imag} */,
  {32'hc2db8334, 32'hc162fde9} /* (6, 5, 20) {real, imag} */,
  {32'hc21a8f7a, 32'hc211d19c} /* (6, 5, 19) {real, imag} */,
  {32'hc0a62b98, 32'h41cadac8} /* (6, 5, 18) {real, imag} */,
  {32'hc1b1462b, 32'hc2472edc} /* (6, 5, 17) {real, imag} */,
  {32'hc22daaf6, 32'h00000000} /* (6, 5, 16) {real, imag} */,
  {32'hc1b1462b, 32'h42472edc} /* (6, 5, 15) {real, imag} */,
  {32'hc0a62b98, 32'hc1cadac8} /* (6, 5, 14) {real, imag} */,
  {32'hc21a8f7a, 32'h4211d19c} /* (6, 5, 13) {real, imag} */,
  {32'hc2db8334, 32'h4162fde9} /* (6, 5, 12) {real, imag} */,
  {32'hc2b7f392, 32'hc2859a0b} /* (6, 5, 11) {real, imag} */,
  {32'h43131105, 32'h422bd33b} /* (6, 5, 10) {real, imag} */,
  {32'hc2d084f6, 32'h42f1d38e} /* (6, 5, 9) {real, imag} */,
  {32'hc09ddfb8, 32'h417d5c52} /* (6, 5, 8) {real, imag} */,
  {32'h42869de8, 32'h429d56c4} /* (6, 5, 7) {real, imag} */,
  {32'h425e7127, 32'h40bc862c} /* (6, 5, 6) {real, imag} */,
  {32'hc2ec9173, 32'h42b9705b} /* (6, 5, 5) {real, imag} */,
  {32'h41cab508, 32'hc095f160} /* (6, 5, 4) {real, imag} */,
  {32'h41e28a5c, 32'hc26a9ae3} /* (6, 5, 3) {real, imag} */,
  {32'hc31cc9c4, 32'hc420e3ca} /* (6, 5, 2) {real, imag} */,
  {32'h44efa338, 32'h44c32180} /* (6, 5, 1) {real, imag} */,
  {32'h453960f3, 32'h00000000} /* (6, 5, 0) {real, imag} */,
  {32'h44e797b9, 32'hc4ef8c0e} /* (6, 4, 31) {real, imag} */,
  {32'h4311671c, 32'h4447635e} /* (6, 4, 30) {real, imag} */,
  {32'h4315e27c, 32'h41be36eb} /* (6, 4, 29) {real, imag} */,
  {32'hc291d121, 32'h43a4d910} /* (6, 4, 28) {real, imag} */,
  {32'hc244f00c, 32'hc2e5122e} /* (6, 4, 27) {real, imag} */,
  {32'h4289ca14, 32'h42508fce} /* (6, 4, 26) {real, imag} */,
  {32'h42d563ca, 32'hc2e4eccc} /* (6, 4, 25) {real, imag} */,
  {32'h4281a9bb, 32'h42e454c2} /* (6, 4, 24) {real, imag} */,
  {32'hc25feae2, 32'hc1fe2db0} /* (6, 4, 23) {real, imag} */,
  {32'h42a7be20, 32'h42dc00df} /* (6, 4, 22) {real, imag} */,
  {32'hc26fa3da, 32'h40548800} /* (6, 4, 21) {real, imag} */,
  {32'hc2271fc8, 32'h41a57453} /* (6, 4, 20) {real, imag} */,
  {32'hc2d64344, 32'h4253c715} /* (6, 4, 19) {real, imag} */,
  {32'hc1856f68, 32'hc255b45e} /* (6, 4, 18) {real, imag} */,
  {32'hc2a20b00, 32'h42d76f4d} /* (6, 4, 17) {real, imag} */,
  {32'h416411e2, 32'h00000000} /* (6, 4, 16) {real, imag} */,
  {32'hc2a20b00, 32'hc2d76f4d} /* (6, 4, 15) {real, imag} */,
  {32'hc1856f68, 32'h4255b45e} /* (6, 4, 14) {real, imag} */,
  {32'hc2d64344, 32'hc253c715} /* (6, 4, 13) {real, imag} */,
  {32'hc2271fc8, 32'hc1a57453} /* (6, 4, 12) {real, imag} */,
  {32'hc26fa3da, 32'hc0548800} /* (6, 4, 11) {real, imag} */,
  {32'h42a7be20, 32'hc2dc00df} /* (6, 4, 10) {real, imag} */,
  {32'hc25feae2, 32'h41fe2db0} /* (6, 4, 9) {real, imag} */,
  {32'h4281a9bb, 32'hc2e454c2} /* (6, 4, 8) {real, imag} */,
  {32'h42d563ca, 32'h42e4eccc} /* (6, 4, 7) {real, imag} */,
  {32'h4289ca14, 32'hc2508fce} /* (6, 4, 6) {real, imag} */,
  {32'hc244f00c, 32'h42e5122e} /* (6, 4, 5) {real, imag} */,
  {32'hc291d121, 32'hc3a4d910} /* (6, 4, 4) {real, imag} */,
  {32'h4315e27c, 32'hc1be36eb} /* (6, 4, 3) {real, imag} */,
  {32'h4311671c, 32'hc447635e} /* (6, 4, 2) {real, imag} */,
  {32'h44e797b9, 32'h44ef8c0e} /* (6, 4, 1) {real, imag} */,
  {32'h453ada56, 32'h00000000} /* (6, 4, 0) {real, imag} */,
  {32'h44da23ce, 32'hc5027e74} /* (6, 3, 31) {real, imag} */,
  {32'h433cf5da, 32'h4419ee10} /* (6, 3, 30) {real, imag} */,
  {32'h41f2a142, 32'h42174284} /* (6, 3, 29) {real, imag} */,
  {32'h41e1c178, 32'h434ded56} /* (6, 3, 28) {real, imag} */,
  {32'hc29c32e5, 32'hc2c17e00} /* (6, 3, 27) {real, imag} */,
  {32'h40b885c8, 32'h4199489b} /* (6, 3, 26) {real, imag} */,
  {32'h41f1f503, 32'hc232c329} /* (6, 3, 25) {real, imag} */,
  {32'h42de13dd, 32'h41c80881} /* (6, 3, 24) {real, imag} */,
  {32'h4297fc97, 32'hc09ccb08} /* (6, 3, 23) {real, imag} */,
  {32'h41932661, 32'h41c6eda1} /* (6, 3, 22) {real, imag} */,
  {32'hc2fc0188, 32'h42d42c55} /* (6, 3, 21) {real, imag} */,
  {32'h4084cf26, 32'hc0e3e79c} /* (6, 3, 20) {real, imag} */,
  {32'h4235b681, 32'h42a6d838} /* (6, 3, 19) {real, imag} */,
  {32'hc246e581, 32'h40811630} /* (6, 3, 18) {real, imag} */,
  {32'h41eab584, 32'h4201b1ce} /* (6, 3, 17) {real, imag} */,
  {32'hc17b62d6, 32'h00000000} /* (6, 3, 16) {real, imag} */,
  {32'h41eab584, 32'hc201b1ce} /* (6, 3, 15) {real, imag} */,
  {32'hc246e581, 32'hc0811630} /* (6, 3, 14) {real, imag} */,
  {32'h4235b681, 32'hc2a6d838} /* (6, 3, 13) {real, imag} */,
  {32'h4084cf26, 32'h40e3e79c} /* (6, 3, 12) {real, imag} */,
  {32'hc2fc0188, 32'hc2d42c55} /* (6, 3, 11) {real, imag} */,
  {32'h41932661, 32'hc1c6eda1} /* (6, 3, 10) {real, imag} */,
  {32'h4297fc97, 32'h409ccb08} /* (6, 3, 9) {real, imag} */,
  {32'h42de13dd, 32'hc1c80881} /* (6, 3, 8) {real, imag} */,
  {32'h41f1f503, 32'h4232c329} /* (6, 3, 7) {real, imag} */,
  {32'h40b885c8, 32'hc199489b} /* (6, 3, 6) {real, imag} */,
  {32'hc29c32e5, 32'h42c17e00} /* (6, 3, 5) {real, imag} */,
  {32'h41e1c178, 32'hc34ded56} /* (6, 3, 4) {real, imag} */,
  {32'h41f2a142, 32'hc2174284} /* (6, 3, 3) {real, imag} */,
  {32'h433cf5da, 32'hc419ee10} /* (6, 3, 2) {real, imag} */,
  {32'h44da23ce, 32'h45027e74} /* (6, 3, 1) {real, imag} */,
  {32'h4549922c, 32'h00000000} /* (6, 3, 0) {real, imag} */,
  {32'h44c70934, 32'hc503bb85} /* (6, 2, 31) {real, imag} */,
  {32'h435abc1c, 32'h44127cd2} /* (6, 2, 30) {real, imag} */,
  {32'h4200d836, 32'h42241df4} /* (6, 2, 29) {real, imag} */,
  {32'h419bfb3a, 32'h42cec554} /* (6, 2, 28) {real, imag} */,
  {32'hc30dad0c, 32'hc0b83828} /* (6, 2, 27) {real, imag} */,
  {32'h410132c3, 32'h426af036} /* (6, 2, 26) {real, imag} */,
  {32'hc1e08e34, 32'hc2809b41} /* (6, 2, 25) {real, imag} */,
  {32'h41ae1a3b, 32'h42e4649b} /* (6, 2, 24) {real, imag} */,
  {32'hc23139ed, 32'hc2aaa7c9} /* (6, 2, 23) {real, imag} */,
  {32'hc11dacfc, 32'hc3045306} /* (6, 2, 22) {real, imag} */,
  {32'hc2a0cd47, 32'h40850930} /* (6, 2, 21) {real, imag} */,
  {32'h4248e245, 32'h42fdaf0e} /* (6, 2, 20) {real, imag} */,
  {32'h42e1f2c8, 32'hc14a33a0} /* (6, 2, 19) {real, imag} */,
  {32'h42467317, 32'hc21f62ff} /* (6, 2, 18) {real, imag} */,
  {32'h42379bfc, 32'h429a7532} /* (6, 2, 17) {real, imag} */,
  {32'h4207ee52, 32'h00000000} /* (6, 2, 16) {real, imag} */,
  {32'h42379bfc, 32'hc29a7532} /* (6, 2, 15) {real, imag} */,
  {32'h42467317, 32'h421f62ff} /* (6, 2, 14) {real, imag} */,
  {32'h42e1f2c8, 32'h414a33a0} /* (6, 2, 13) {real, imag} */,
  {32'h4248e245, 32'hc2fdaf0e} /* (6, 2, 12) {real, imag} */,
  {32'hc2a0cd47, 32'hc0850930} /* (6, 2, 11) {real, imag} */,
  {32'hc11dacfc, 32'h43045306} /* (6, 2, 10) {real, imag} */,
  {32'hc23139ed, 32'h42aaa7c9} /* (6, 2, 9) {real, imag} */,
  {32'h41ae1a3b, 32'hc2e4649b} /* (6, 2, 8) {real, imag} */,
  {32'hc1e08e34, 32'h42809b41} /* (6, 2, 7) {real, imag} */,
  {32'h410132c3, 32'hc26af036} /* (6, 2, 6) {real, imag} */,
  {32'hc30dad0c, 32'h40b83828} /* (6, 2, 5) {real, imag} */,
  {32'h419bfb3a, 32'hc2cec554} /* (6, 2, 4) {real, imag} */,
  {32'h4200d836, 32'hc2241df4} /* (6, 2, 3) {real, imag} */,
  {32'h435abc1c, 32'hc4127cd2} /* (6, 2, 2) {real, imag} */,
  {32'h44c70934, 32'h4503bb85} /* (6, 2, 1) {real, imag} */,
  {32'h4566f35f, 32'h00000000} /* (6, 2, 0) {real, imag} */,
  {32'h44ce42cf, 32'hc4e521ce} /* (6, 1, 31) {real, imag} */,
  {32'h43395200, 32'h43c38656} /* (6, 1, 30) {real, imag} */,
  {32'hc2d6e5a6, 32'h42499c56} /* (6, 1, 29) {real, imag} */,
  {32'hc07b6410, 32'h42584265} /* (6, 1, 28) {real, imag} */,
  {32'hc2cd6ed6, 32'h41dbf5bf} /* (6, 1, 27) {real, imag} */,
  {32'hc107f280, 32'hc0dbc8bc} /* (6, 1, 26) {real, imag} */,
  {32'h424d197e, 32'hc23c86c3} /* (6, 1, 25) {real, imag} */,
  {32'hc187042b, 32'h42a1e0d1} /* (6, 1, 24) {real, imag} */,
  {32'h423b410f, 32'hc2133930} /* (6, 1, 23) {real, imag} */,
  {32'hc27de8bb, 32'hc05480e0} /* (6, 1, 22) {real, imag} */,
  {32'h41bfa981, 32'h40f3352c} /* (6, 1, 21) {real, imag} */,
  {32'hc19e6778, 32'h418f895d} /* (6, 1, 20) {real, imag} */,
  {32'h421a9cb6, 32'h4192eff2} /* (6, 1, 19) {real, imag} */,
  {32'h41e9c4bd, 32'h421f7032} /* (6, 1, 18) {real, imag} */,
  {32'hc2ae9402, 32'h4047a636} /* (6, 1, 17) {real, imag} */,
  {32'hc1b48955, 32'h00000000} /* (6, 1, 16) {real, imag} */,
  {32'hc2ae9402, 32'hc047a636} /* (6, 1, 15) {real, imag} */,
  {32'h41e9c4bd, 32'hc21f7032} /* (6, 1, 14) {real, imag} */,
  {32'h421a9cb6, 32'hc192eff2} /* (6, 1, 13) {real, imag} */,
  {32'hc19e6778, 32'hc18f895d} /* (6, 1, 12) {real, imag} */,
  {32'h41bfa981, 32'hc0f3352c} /* (6, 1, 11) {real, imag} */,
  {32'hc27de8bb, 32'h405480e0} /* (6, 1, 10) {real, imag} */,
  {32'h423b410f, 32'h42133930} /* (6, 1, 9) {real, imag} */,
  {32'hc187042b, 32'hc2a1e0d1} /* (6, 1, 8) {real, imag} */,
  {32'h424d197e, 32'h423c86c3} /* (6, 1, 7) {real, imag} */,
  {32'hc107f280, 32'h40dbc8bc} /* (6, 1, 6) {real, imag} */,
  {32'hc2cd6ed6, 32'hc1dbf5bf} /* (6, 1, 5) {real, imag} */,
  {32'hc07b6410, 32'hc2584265} /* (6, 1, 4) {real, imag} */,
  {32'hc2d6e5a6, 32'hc2499c56} /* (6, 1, 3) {real, imag} */,
  {32'h43395200, 32'hc3c38656} /* (6, 1, 2) {real, imag} */,
  {32'h44ce42cf, 32'h44e521ce} /* (6, 1, 1) {real, imag} */,
  {32'h455828e7, 32'h00000000} /* (6, 1, 0) {real, imag} */,
  {32'h44e83bf9, 32'hc4bc41a5} /* (6, 0, 31) {real, imag} */,
  {32'hc137a1a0, 32'h438d1cb4} /* (6, 0, 30) {real, imag} */,
  {32'hc29c1b6b, 32'h412090c2} /* (6, 0, 29) {real, imag} */,
  {32'hc2595b27, 32'h4298056a} /* (6, 0, 28) {real, imag} */,
  {32'hc25edc13, 32'h42064ccd} /* (6, 0, 27) {real, imag} */,
  {32'h42445293, 32'hc2c82ae4} /* (6, 0, 26) {real, imag} */,
  {32'h42404f68, 32'hc264fc60} /* (6, 0, 25) {real, imag} */,
  {32'hc0394200, 32'hc197a4d0} /* (6, 0, 24) {real, imag} */,
  {32'hc04cf6f8, 32'hc28db562} /* (6, 0, 23) {real, imag} */,
  {32'hc2e0770e, 32'h42778b18} /* (6, 0, 22) {real, imag} */,
  {32'hc1e326a6, 32'h41c6ae84} /* (6, 0, 21) {real, imag} */,
  {32'h423cc262, 32'h41d50c1d} /* (6, 0, 20) {real, imag} */,
  {32'h4208e99a, 32'hc0d06a68} /* (6, 0, 19) {real, imag} */,
  {32'h425adc58, 32'hc256952e} /* (6, 0, 18) {real, imag} */,
  {32'hc25a8976, 32'hc28171be} /* (6, 0, 17) {real, imag} */,
  {32'hc288ab5e, 32'h00000000} /* (6, 0, 16) {real, imag} */,
  {32'hc25a8976, 32'h428171be} /* (6, 0, 15) {real, imag} */,
  {32'h425adc58, 32'h4256952e} /* (6, 0, 14) {real, imag} */,
  {32'h4208e99a, 32'h40d06a68} /* (6, 0, 13) {real, imag} */,
  {32'h423cc262, 32'hc1d50c1d} /* (6, 0, 12) {real, imag} */,
  {32'hc1e326a6, 32'hc1c6ae84} /* (6, 0, 11) {real, imag} */,
  {32'hc2e0770e, 32'hc2778b18} /* (6, 0, 10) {real, imag} */,
  {32'hc04cf6f8, 32'h428db562} /* (6, 0, 9) {real, imag} */,
  {32'hc0394200, 32'h4197a4d0} /* (6, 0, 8) {real, imag} */,
  {32'h42404f68, 32'h4264fc60} /* (6, 0, 7) {real, imag} */,
  {32'h42445293, 32'h42c82ae4} /* (6, 0, 6) {real, imag} */,
  {32'hc25edc13, 32'hc2064ccd} /* (6, 0, 5) {real, imag} */,
  {32'hc2595b27, 32'hc298056a} /* (6, 0, 4) {real, imag} */,
  {32'hc29c1b6b, 32'hc12090c2} /* (6, 0, 3) {real, imag} */,
  {32'hc137a1a0, 32'hc38d1cb4} /* (6, 0, 2) {real, imag} */,
  {32'h44e83bf9, 32'h44bc41a5} /* (6, 0, 1) {real, imag} */,
  {32'h45554f8c, 32'h00000000} /* (6, 0, 0) {real, imag} */,
  {32'h445d5fd4, 32'hc40542d1} /* (5, 31, 31) {real, imag} */,
  {32'h41a0a4ff, 32'hc2b8b24b} /* (5, 31, 30) {real, imag} */,
  {32'h42b15579, 32'hc2ccf1d7} /* (5, 31, 29) {real, imag} */,
  {32'h41fbc713, 32'hc1eba626} /* (5, 31, 28) {real, imag} */,
  {32'h4227ce59, 32'hc1dabb75} /* (5, 31, 27) {real, imag} */,
  {32'h428266b9, 32'h42189215} /* (5, 31, 26) {real, imag} */,
  {32'h40caabcc, 32'h4223ed12} /* (5, 31, 25) {real, imag} */,
  {32'hc05345c0, 32'h42142070} /* (5, 31, 24) {real, imag} */,
  {32'h4205e63e, 32'h420c22d7} /* (5, 31, 23) {real, imag} */,
  {32'h403e5e1c, 32'hc1cff522} /* (5, 31, 22) {real, imag} */,
  {32'hc27d151b, 32'h42a2aefd} /* (5, 31, 21) {real, imag} */,
  {32'h40b43f30, 32'hc2350372} /* (5, 31, 20) {real, imag} */,
  {32'h41131f70, 32'h42547f60} /* (5, 31, 19) {real, imag} */,
  {32'h413e3374, 32'hc11ae4b0} /* (5, 31, 18) {real, imag} */,
  {32'h419534da, 32'hc16c3a92} /* (5, 31, 17) {real, imag} */,
  {32'hc20dbd9e, 32'h00000000} /* (5, 31, 16) {real, imag} */,
  {32'h419534da, 32'h416c3a92} /* (5, 31, 15) {real, imag} */,
  {32'h413e3374, 32'h411ae4b0} /* (5, 31, 14) {real, imag} */,
  {32'h41131f70, 32'hc2547f60} /* (5, 31, 13) {real, imag} */,
  {32'h40b43f30, 32'h42350372} /* (5, 31, 12) {real, imag} */,
  {32'hc27d151b, 32'hc2a2aefd} /* (5, 31, 11) {real, imag} */,
  {32'h403e5e1c, 32'h41cff522} /* (5, 31, 10) {real, imag} */,
  {32'h4205e63e, 32'hc20c22d7} /* (5, 31, 9) {real, imag} */,
  {32'hc05345c0, 32'hc2142070} /* (5, 31, 8) {real, imag} */,
  {32'h40caabcc, 32'hc223ed12} /* (5, 31, 7) {real, imag} */,
  {32'h428266b9, 32'hc2189215} /* (5, 31, 6) {real, imag} */,
  {32'h4227ce59, 32'h41dabb75} /* (5, 31, 5) {real, imag} */,
  {32'h41fbc713, 32'h41eba626} /* (5, 31, 4) {real, imag} */,
  {32'h42b15579, 32'h42ccf1d7} /* (5, 31, 3) {real, imag} */,
  {32'h41a0a4ff, 32'h42b8b24b} /* (5, 31, 2) {real, imag} */,
  {32'h445d5fd4, 32'h440542d1} /* (5, 31, 1) {real, imag} */,
  {32'h450035c1, 32'h00000000} /* (5, 31, 0) {real, imag} */,
  {32'h445d21d9, 32'hc3f9f656} /* (5, 30, 31) {real, imag} */,
  {32'h4335598c, 32'hc2730125} /* (5, 30, 30) {real, imag} */,
  {32'h4325aaab, 32'hc2df0ab6} /* (5, 30, 29) {real, imag} */,
  {32'h42804c35, 32'h41e3f558} /* (5, 30, 28) {real, imag} */,
  {32'hc21efd91, 32'h42b268f6} /* (5, 30, 27) {real, imag} */,
  {32'hc24c4d2a, 32'h4292a631} /* (5, 30, 26) {real, imag} */,
  {32'hc30d0dd1, 32'hc12cee08} /* (5, 30, 25) {real, imag} */,
  {32'h42cd7b9d, 32'hc23d1f59} /* (5, 30, 24) {real, imag} */,
  {32'h41f69ad8, 32'hc24b4842} /* (5, 30, 23) {real, imag} */,
  {32'hc2aabe3d, 32'h4308fb2d} /* (5, 30, 22) {real, imag} */,
  {32'h4250d849, 32'h4292a57b} /* (5, 30, 21) {real, imag} */,
  {32'hc10ca4ca, 32'hc262c336} /* (5, 30, 20) {real, imag} */,
  {32'h4226b186, 32'hc04abd88} /* (5, 30, 19) {real, imag} */,
  {32'h4242f6d2, 32'h41bf35d3} /* (5, 30, 18) {real, imag} */,
  {32'h416342a1, 32'hc1aa38ec} /* (5, 30, 17) {real, imag} */,
  {32'hc2846469, 32'h00000000} /* (5, 30, 16) {real, imag} */,
  {32'h416342a1, 32'h41aa38ec} /* (5, 30, 15) {real, imag} */,
  {32'h4242f6d2, 32'hc1bf35d3} /* (5, 30, 14) {real, imag} */,
  {32'h4226b186, 32'h404abd88} /* (5, 30, 13) {real, imag} */,
  {32'hc10ca4ca, 32'h4262c336} /* (5, 30, 12) {real, imag} */,
  {32'h4250d849, 32'hc292a57b} /* (5, 30, 11) {real, imag} */,
  {32'hc2aabe3d, 32'hc308fb2d} /* (5, 30, 10) {real, imag} */,
  {32'h41f69ad8, 32'h424b4842} /* (5, 30, 9) {real, imag} */,
  {32'h42cd7b9d, 32'h423d1f59} /* (5, 30, 8) {real, imag} */,
  {32'hc30d0dd1, 32'h412cee08} /* (5, 30, 7) {real, imag} */,
  {32'hc24c4d2a, 32'hc292a631} /* (5, 30, 6) {real, imag} */,
  {32'hc21efd91, 32'hc2b268f6} /* (5, 30, 5) {real, imag} */,
  {32'h42804c35, 32'hc1e3f558} /* (5, 30, 4) {real, imag} */,
  {32'h4325aaab, 32'h42df0ab6} /* (5, 30, 3) {real, imag} */,
  {32'h4335598c, 32'h42730125} /* (5, 30, 2) {real, imag} */,
  {32'h445d21d9, 32'h43f9f656} /* (5, 30, 1) {real, imag} */,
  {32'h45040d9a, 32'h00000000} /* (5, 30, 0) {real, imag} */,
  {32'h44516f18, 32'hc38871d0} /* (5, 29, 31) {real, imag} */,
  {32'h433acb88, 32'h423c2968} /* (5, 29, 30) {real, imag} */,
  {32'h431f8669, 32'hc1b02f20} /* (5, 29, 29) {real, imag} */,
  {32'h42cdf156, 32'hc27ac194} /* (5, 29, 28) {real, imag} */,
  {32'hc123d76c, 32'h432156c8} /* (5, 29, 27) {real, imag} */,
  {32'hc1e335cc, 32'h42aa2ffa} /* (5, 29, 26) {real, imag} */,
  {32'hc2182bad, 32'hc2f5db6a} /* (5, 29, 25) {real, imag} */,
  {32'h430a2ef5, 32'hc2cfbc2c} /* (5, 29, 24) {real, imag} */,
  {32'h418cc474, 32'hc29cc018} /* (5, 29, 23) {real, imag} */,
  {32'hc31b1bad, 32'h4047bc40} /* (5, 29, 22) {real, imag} */,
  {32'hc298692c, 32'h40b8db2c} /* (5, 29, 21) {real, imag} */,
  {32'h4214b246, 32'hc0a3fd80} /* (5, 29, 20) {real, imag} */,
  {32'h420dd6a5, 32'h419d9564} /* (5, 29, 19) {real, imag} */,
  {32'hc2242d0f, 32'h4314fc16} /* (5, 29, 18) {real, imag} */,
  {32'h3f7b5820, 32'h42735aef} /* (5, 29, 17) {real, imag} */,
  {32'h4088efec, 32'h00000000} /* (5, 29, 16) {real, imag} */,
  {32'h3f7b5820, 32'hc2735aef} /* (5, 29, 15) {real, imag} */,
  {32'hc2242d0f, 32'hc314fc16} /* (5, 29, 14) {real, imag} */,
  {32'h420dd6a5, 32'hc19d9564} /* (5, 29, 13) {real, imag} */,
  {32'h4214b246, 32'h40a3fd80} /* (5, 29, 12) {real, imag} */,
  {32'hc298692c, 32'hc0b8db2c} /* (5, 29, 11) {real, imag} */,
  {32'hc31b1bad, 32'hc047bc40} /* (5, 29, 10) {real, imag} */,
  {32'h418cc474, 32'h429cc018} /* (5, 29, 9) {real, imag} */,
  {32'h430a2ef5, 32'h42cfbc2c} /* (5, 29, 8) {real, imag} */,
  {32'hc2182bad, 32'h42f5db6a} /* (5, 29, 7) {real, imag} */,
  {32'hc1e335cc, 32'hc2aa2ffa} /* (5, 29, 6) {real, imag} */,
  {32'hc123d76c, 32'hc32156c8} /* (5, 29, 5) {real, imag} */,
  {32'h42cdf156, 32'h427ac194} /* (5, 29, 4) {real, imag} */,
  {32'h431f8669, 32'h41b02f20} /* (5, 29, 3) {real, imag} */,
  {32'h433acb88, 32'hc23c2968} /* (5, 29, 2) {real, imag} */,
  {32'h44516f18, 32'h438871d0} /* (5, 29, 1) {real, imag} */,
  {32'h44ec01a5, 32'h00000000} /* (5, 29, 0) {real, imag} */,
  {32'h442bc93a, 32'hc31148f4} /* (5, 28, 31) {real, imag} */,
  {32'h41eee107, 32'h4181cc34} /* (5, 28, 30) {real, imag} */,
  {32'h435717bf, 32'h41eb83b0} /* (5, 28, 29) {real, imag} */,
  {32'hc2982130, 32'h41c76b33} /* (5, 28, 28) {real, imag} */,
  {32'hc2bae2f4, 32'hc23bd256} /* (5, 28, 27) {real, imag} */,
  {32'h43097ac1, 32'h40431428} /* (5, 28, 26) {real, imag} */,
  {32'h425490b0, 32'h41b1dbf0} /* (5, 28, 25) {real, imag} */,
  {32'h428d2998, 32'h3ff387d0} /* (5, 28, 24) {real, imag} */,
  {32'h424aabb0, 32'hc304f5b3} /* (5, 28, 23) {real, imag} */,
  {32'hc246efe6, 32'hc279a8f0} /* (5, 28, 22) {real, imag} */,
  {32'hc2ac6a20, 32'h42ccb767} /* (5, 28, 21) {real, imag} */,
  {32'hc1eae2c1, 32'hc29624f9} /* (5, 28, 20) {real, imag} */,
  {32'h400b01a8, 32'hc241b43b} /* (5, 28, 19) {real, imag} */,
  {32'hc2a17fea, 32'h4100d870} /* (5, 28, 18) {real, imag} */,
  {32'hc20379f5, 32'hc2703a7f} /* (5, 28, 17) {real, imag} */,
  {32'h4280cf8d, 32'h00000000} /* (5, 28, 16) {real, imag} */,
  {32'hc20379f5, 32'h42703a7f} /* (5, 28, 15) {real, imag} */,
  {32'hc2a17fea, 32'hc100d870} /* (5, 28, 14) {real, imag} */,
  {32'h400b01a8, 32'h4241b43b} /* (5, 28, 13) {real, imag} */,
  {32'hc1eae2c1, 32'h429624f9} /* (5, 28, 12) {real, imag} */,
  {32'hc2ac6a20, 32'hc2ccb767} /* (5, 28, 11) {real, imag} */,
  {32'hc246efe6, 32'h4279a8f0} /* (5, 28, 10) {real, imag} */,
  {32'h424aabb0, 32'h4304f5b3} /* (5, 28, 9) {real, imag} */,
  {32'h428d2998, 32'hbff387d0} /* (5, 28, 8) {real, imag} */,
  {32'h425490b0, 32'hc1b1dbf0} /* (5, 28, 7) {real, imag} */,
  {32'h43097ac1, 32'hc0431428} /* (5, 28, 6) {real, imag} */,
  {32'hc2bae2f4, 32'h423bd256} /* (5, 28, 5) {real, imag} */,
  {32'hc2982130, 32'hc1c76b33} /* (5, 28, 4) {real, imag} */,
  {32'h435717bf, 32'hc1eb83b0} /* (5, 28, 3) {real, imag} */,
  {32'h41eee107, 32'hc181cc34} /* (5, 28, 2) {real, imag} */,
  {32'h442bc93a, 32'h431148f4} /* (5, 28, 1) {real, imag} */,
  {32'h44ecdf92, 32'h00000000} /* (5, 28, 0) {real, imag} */,
  {32'h440aeea5, 32'h422fc694} /* (5, 27, 31) {real, imag} */,
  {32'hc10ec7cc, 32'h426607a4} /* (5, 27, 30) {real, imag} */,
  {32'h431a1748, 32'hc3209dc6} /* (5, 27, 29) {real, imag} */,
  {32'hc2f55f4a, 32'hc1bc1804} /* (5, 27, 28) {real, imag} */,
  {32'hc10ac318, 32'h42248c21} /* (5, 27, 27) {real, imag} */,
  {32'h42e04108, 32'hc1f8242d} /* (5, 27, 26) {real, imag} */,
  {32'hc2d299a6, 32'hc109e8c8} /* (5, 27, 25) {real, imag} */,
  {32'hc228d36f, 32'h420d0964} /* (5, 27, 24) {real, imag} */,
  {32'h41112bfc, 32'h42a0abb3} /* (5, 27, 23) {real, imag} */,
  {32'h4268d25e, 32'hc0b990bc} /* (5, 27, 22) {real, imag} */,
  {32'hc08184b0, 32'hc2a6f3f8} /* (5, 27, 21) {real, imag} */,
  {32'hc23ec31c, 32'hc28ccd15} /* (5, 27, 20) {real, imag} */,
  {32'hc2b4d452, 32'h41becc44} /* (5, 27, 19) {real, imag} */,
  {32'hc2260dca, 32'hc249c4bd} /* (5, 27, 18) {real, imag} */,
  {32'h41b50b3a, 32'hc05b8250} /* (5, 27, 17) {real, imag} */,
  {32'hc2e855b4, 32'h00000000} /* (5, 27, 16) {real, imag} */,
  {32'h41b50b3a, 32'h405b8250} /* (5, 27, 15) {real, imag} */,
  {32'hc2260dca, 32'h4249c4bd} /* (5, 27, 14) {real, imag} */,
  {32'hc2b4d452, 32'hc1becc44} /* (5, 27, 13) {real, imag} */,
  {32'hc23ec31c, 32'h428ccd15} /* (5, 27, 12) {real, imag} */,
  {32'hc08184b0, 32'h42a6f3f8} /* (5, 27, 11) {real, imag} */,
  {32'h4268d25e, 32'h40b990bc} /* (5, 27, 10) {real, imag} */,
  {32'h41112bfc, 32'hc2a0abb3} /* (5, 27, 9) {real, imag} */,
  {32'hc228d36f, 32'hc20d0964} /* (5, 27, 8) {real, imag} */,
  {32'hc2d299a6, 32'h4109e8c8} /* (5, 27, 7) {real, imag} */,
  {32'h42e04108, 32'h41f8242d} /* (5, 27, 6) {real, imag} */,
  {32'hc10ac318, 32'hc2248c21} /* (5, 27, 5) {real, imag} */,
  {32'hc2f55f4a, 32'h41bc1804} /* (5, 27, 4) {real, imag} */,
  {32'h431a1748, 32'h43209dc6} /* (5, 27, 3) {real, imag} */,
  {32'hc10ec7cc, 32'hc26607a4} /* (5, 27, 2) {real, imag} */,
  {32'h440aeea5, 32'hc22fc694} /* (5, 27, 1) {real, imag} */,
  {32'h44e23158, 32'h00000000} /* (5, 27, 0) {real, imag} */,
  {32'h440edde5, 32'h4100ea90} /* (5, 26, 31) {real, imag} */,
  {32'h41df155a, 32'h4296c0f8} /* (5, 26, 30) {real, imag} */,
  {32'hc2329850, 32'hc30f2679} /* (5, 26, 29) {real, imag} */,
  {32'hc22634c2, 32'hc0af81a0} /* (5, 26, 28) {real, imag} */,
  {32'h42a36620, 32'h42d342a2} /* (5, 26, 27) {real, imag} */,
  {32'hc1551341, 32'hc1932b1d} /* (5, 26, 26) {real, imag} */,
  {32'hc0f2cc7c, 32'hc25a238c} /* (5, 26, 25) {real, imag} */,
  {32'hc298e7e2, 32'hc28001c5} /* (5, 26, 24) {real, imag} */,
  {32'hc2229b3e, 32'h430b5586} /* (5, 26, 23) {real, imag} */,
  {32'hc28b51ab, 32'hc1cfdfdc} /* (5, 26, 22) {real, imag} */,
  {32'h4256eae6, 32'h41ca1476} /* (5, 26, 21) {real, imag} */,
  {32'hc2c03bc2, 32'h408e9d20} /* (5, 26, 20) {real, imag} */,
  {32'hc1aeb0df, 32'h41830854} /* (5, 26, 19) {real, imag} */,
  {32'hbfd7bb00, 32'hc1bee2e3} /* (5, 26, 18) {real, imag} */,
  {32'hc1e4f5c0, 32'hbfefbd78} /* (5, 26, 17) {real, imag} */,
  {32'h4271ffec, 32'h00000000} /* (5, 26, 16) {real, imag} */,
  {32'hc1e4f5c0, 32'h3fefbd78} /* (5, 26, 15) {real, imag} */,
  {32'hbfd7bb00, 32'h41bee2e3} /* (5, 26, 14) {real, imag} */,
  {32'hc1aeb0df, 32'hc1830854} /* (5, 26, 13) {real, imag} */,
  {32'hc2c03bc2, 32'hc08e9d20} /* (5, 26, 12) {real, imag} */,
  {32'h4256eae6, 32'hc1ca1476} /* (5, 26, 11) {real, imag} */,
  {32'hc28b51ab, 32'h41cfdfdc} /* (5, 26, 10) {real, imag} */,
  {32'hc2229b3e, 32'hc30b5586} /* (5, 26, 9) {real, imag} */,
  {32'hc298e7e2, 32'h428001c5} /* (5, 26, 8) {real, imag} */,
  {32'hc0f2cc7c, 32'h425a238c} /* (5, 26, 7) {real, imag} */,
  {32'hc1551341, 32'h41932b1d} /* (5, 26, 6) {real, imag} */,
  {32'h42a36620, 32'hc2d342a2} /* (5, 26, 5) {real, imag} */,
  {32'hc22634c2, 32'h40af81a0} /* (5, 26, 4) {real, imag} */,
  {32'hc2329850, 32'h430f2679} /* (5, 26, 3) {real, imag} */,
  {32'h41df155a, 32'hc296c0f8} /* (5, 26, 2) {real, imag} */,
  {32'h440edde5, 32'hc100ea90} /* (5, 26, 1) {real, imag} */,
  {32'h44dcc66c, 32'h00000000} /* (5, 26, 0) {real, imag} */,
  {32'h439266f6, 32'hc0a89f20} /* (5, 25, 31) {real, imag} */,
  {32'h429fa41c, 32'h42a68e40} /* (5, 25, 30) {real, imag} */,
  {32'hc2b86666, 32'hc2f5fbe1} /* (5, 25, 29) {real, imag} */,
  {32'hc2bff5b6, 32'h411d2ee4} /* (5, 25, 28) {real, imag} */,
  {32'h42d170c6, 32'hc216cdc4} /* (5, 25, 27) {real, imag} */,
  {32'h431be93c, 32'hc20f2186} /* (5, 25, 26) {real, imag} */,
  {32'h42a7f70f, 32'h42b0e4bc} /* (5, 25, 25) {real, imag} */,
  {32'h418591f1, 32'hc1ec2308} /* (5, 25, 24) {real, imag} */,
  {32'hc1d1a208, 32'h41fb1f7e} /* (5, 25, 23) {real, imag} */,
  {32'hc1b08bda, 32'h4203d854} /* (5, 25, 22) {real, imag} */,
  {32'h427e554a, 32'hc275bcb6} /* (5, 25, 21) {real, imag} */,
  {32'hc3109f66, 32'h429a05f8} /* (5, 25, 20) {real, imag} */,
  {32'h4209010a, 32'hc23d2028} /* (5, 25, 19) {real, imag} */,
  {32'hc1bb9aa4, 32'hc03df130} /* (5, 25, 18) {real, imag} */,
  {32'hc25e73ab, 32'hc0cb92e8} /* (5, 25, 17) {real, imag} */,
  {32'hc2a4c52c, 32'h00000000} /* (5, 25, 16) {real, imag} */,
  {32'hc25e73ab, 32'h40cb92e8} /* (5, 25, 15) {real, imag} */,
  {32'hc1bb9aa4, 32'h403df130} /* (5, 25, 14) {real, imag} */,
  {32'h4209010a, 32'h423d2028} /* (5, 25, 13) {real, imag} */,
  {32'hc3109f66, 32'hc29a05f8} /* (5, 25, 12) {real, imag} */,
  {32'h427e554a, 32'h4275bcb6} /* (5, 25, 11) {real, imag} */,
  {32'hc1b08bda, 32'hc203d854} /* (5, 25, 10) {real, imag} */,
  {32'hc1d1a208, 32'hc1fb1f7e} /* (5, 25, 9) {real, imag} */,
  {32'h418591f1, 32'h41ec2308} /* (5, 25, 8) {real, imag} */,
  {32'h42a7f70f, 32'hc2b0e4bc} /* (5, 25, 7) {real, imag} */,
  {32'h431be93c, 32'h420f2186} /* (5, 25, 6) {real, imag} */,
  {32'h42d170c6, 32'h4216cdc4} /* (5, 25, 5) {real, imag} */,
  {32'hc2bff5b6, 32'hc11d2ee4} /* (5, 25, 4) {real, imag} */,
  {32'hc2b86666, 32'h42f5fbe1} /* (5, 25, 3) {real, imag} */,
  {32'h429fa41c, 32'hc2a68e40} /* (5, 25, 2) {real, imag} */,
  {32'h439266f6, 32'h40a89f20} /* (5, 25, 1) {real, imag} */,
  {32'h44c13279, 32'h00000000} /* (5, 25, 0) {real, imag} */,
  {32'h4342172f, 32'hc295cb1c} /* (5, 24, 31) {real, imag} */,
  {32'h41a46d98, 32'h430b0fa6} /* (5, 24, 30) {real, imag} */,
  {32'h42b89581, 32'hc30244f8} /* (5, 24, 29) {real, imag} */,
  {32'hc2b6bdee, 32'h40d44570} /* (5, 24, 28) {real, imag} */,
  {32'h42819985, 32'hc303eb5f} /* (5, 24, 27) {real, imag} */,
  {32'h42aebd22, 32'hc2757f84} /* (5, 24, 26) {real, imag} */,
  {32'hc255349e, 32'h42cfd253} /* (5, 24, 25) {real, imag} */,
  {32'h41ef22ca, 32'hc1b2d156} /* (5, 24, 24) {real, imag} */,
  {32'h41fae572, 32'hbf827460} /* (5, 24, 23) {real, imag} */,
  {32'h4230df3c, 32'h42b0b326} /* (5, 24, 22) {real, imag} */,
  {32'hc26e475a, 32'h422574f6} /* (5, 24, 21) {real, imag} */,
  {32'h3f2d7d70, 32'h421b85f0} /* (5, 24, 20) {real, imag} */,
  {32'hc29c148e, 32'h43106fb2} /* (5, 24, 19) {real, imag} */,
  {32'hc233c82b, 32'h42300aee} /* (5, 24, 18) {real, imag} */,
  {32'h419ce4c8, 32'h424aecce} /* (5, 24, 17) {real, imag} */,
  {32'hc26bbb43, 32'h00000000} /* (5, 24, 16) {real, imag} */,
  {32'h419ce4c8, 32'hc24aecce} /* (5, 24, 15) {real, imag} */,
  {32'hc233c82b, 32'hc2300aee} /* (5, 24, 14) {real, imag} */,
  {32'hc29c148e, 32'hc3106fb2} /* (5, 24, 13) {real, imag} */,
  {32'h3f2d7d70, 32'hc21b85f0} /* (5, 24, 12) {real, imag} */,
  {32'hc26e475a, 32'hc22574f6} /* (5, 24, 11) {real, imag} */,
  {32'h4230df3c, 32'hc2b0b326} /* (5, 24, 10) {real, imag} */,
  {32'h41fae572, 32'h3f827460} /* (5, 24, 9) {real, imag} */,
  {32'h41ef22ca, 32'h41b2d156} /* (5, 24, 8) {real, imag} */,
  {32'hc255349e, 32'hc2cfd253} /* (5, 24, 7) {real, imag} */,
  {32'h42aebd22, 32'h42757f84} /* (5, 24, 6) {real, imag} */,
  {32'h42819985, 32'h4303eb5f} /* (5, 24, 5) {real, imag} */,
  {32'hc2b6bdee, 32'hc0d44570} /* (5, 24, 4) {real, imag} */,
  {32'h42b89581, 32'h430244f8} /* (5, 24, 3) {real, imag} */,
  {32'h41a46d98, 32'hc30b0fa6} /* (5, 24, 2) {real, imag} */,
  {32'h4342172f, 32'h4295cb1c} /* (5, 24, 1) {real, imag} */,
  {32'h44af36ff, 32'h00000000} /* (5, 24, 0) {real, imag} */,
  {32'hc21df27a, 32'hc3618b36} /* (5, 23, 31) {real, imag} */,
  {32'h42908105, 32'h423ad840} /* (5, 23, 30) {real, imag} */,
  {32'hc21c66f6, 32'hc2e9342c} /* (5, 23, 29) {real, imag} */,
  {32'hc1b2375b, 32'hc12deeca} /* (5, 23, 28) {real, imag} */,
  {32'h423a80f0, 32'hc2eb029a} /* (5, 23, 27) {real, imag} */,
  {32'hc21ee254, 32'hc2996990} /* (5, 23, 26) {real, imag} */,
  {32'hc2050f32, 32'h411a8fdc} /* (5, 23, 25) {real, imag} */,
  {32'h41c67478, 32'h41d69d1a} /* (5, 23, 24) {real, imag} */,
  {32'h426eea66, 32'hc182bfa2} /* (5, 23, 23) {real, imag} */,
  {32'hc29f3565, 32'h41907c17} /* (5, 23, 22) {real, imag} */,
  {32'h4093d656, 32'h42b089ff} /* (5, 23, 21) {real, imag} */,
  {32'hc1852d9c, 32'h40d45f80} /* (5, 23, 20) {real, imag} */,
  {32'hc149537c, 32'h41bc4f07} /* (5, 23, 19) {real, imag} */,
  {32'hc11d0e4c, 32'h428f97ff} /* (5, 23, 18) {real, imag} */,
  {32'h422dc1cd, 32'hc1d73280} /* (5, 23, 17) {real, imag} */,
  {32'h41bc4300, 32'h00000000} /* (5, 23, 16) {real, imag} */,
  {32'h422dc1cd, 32'h41d73280} /* (5, 23, 15) {real, imag} */,
  {32'hc11d0e4c, 32'hc28f97ff} /* (5, 23, 14) {real, imag} */,
  {32'hc149537c, 32'hc1bc4f07} /* (5, 23, 13) {real, imag} */,
  {32'hc1852d9c, 32'hc0d45f80} /* (5, 23, 12) {real, imag} */,
  {32'h4093d656, 32'hc2b089ff} /* (5, 23, 11) {real, imag} */,
  {32'hc29f3565, 32'hc1907c17} /* (5, 23, 10) {real, imag} */,
  {32'h426eea66, 32'h4182bfa2} /* (5, 23, 9) {real, imag} */,
  {32'h41c67478, 32'hc1d69d1a} /* (5, 23, 8) {real, imag} */,
  {32'hc2050f32, 32'hc11a8fdc} /* (5, 23, 7) {real, imag} */,
  {32'hc21ee254, 32'h42996990} /* (5, 23, 6) {real, imag} */,
  {32'h423a80f0, 32'h42eb029a} /* (5, 23, 5) {real, imag} */,
  {32'hc1b2375b, 32'h412deeca} /* (5, 23, 4) {real, imag} */,
  {32'hc21c66f6, 32'h42e9342c} /* (5, 23, 3) {real, imag} */,
  {32'h42908105, 32'hc23ad840} /* (5, 23, 2) {real, imag} */,
  {32'hc21df27a, 32'h43618b36} /* (5, 23, 1) {real, imag} */,
  {32'h449275e4, 32'h00000000} /* (5, 23, 0) {real, imag} */,
  {32'hc3157118, 32'hc371c773} /* (5, 22, 31) {real, imag} */,
  {32'h41832f84, 32'h42aa38aa} /* (5, 22, 30) {real, imag} */,
  {32'hc281430e, 32'hc33a8b4c} /* (5, 22, 29) {real, imag} */,
  {32'hc2b581d6, 32'h42acd972} /* (5, 22, 28) {real, imag} */,
  {32'h42dc38f9, 32'hc29315aa} /* (5, 22, 27) {real, imag} */,
  {32'h4167edcf, 32'hc22c8b1a} /* (5, 22, 26) {real, imag} */,
  {32'h42775e6e, 32'h4103d9a6} /* (5, 22, 25) {real, imag} */,
  {32'hc1ee2d62, 32'hc25128e4} /* (5, 22, 24) {real, imag} */,
  {32'hc1d997e7, 32'h42a36408} /* (5, 22, 23) {real, imag} */,
  {32'h4232b976, 32'h423d4d03} /* (5, 22, 22) {real, imag} */,
  {32'hc272eea5, 32'h42084db8} /* (5, 22, 21) {real, imag} */,
  {32'hc02f04c0, 32'hc12f7f18} /* (5, 22, 20) {real, imag} */,
  {32'hbfe0ecb0, 32'h41c617f6} /* (5, 22, 19) {real, imag} */,
  {32'h4278778a, 32'hc2328223} /* (5, 22, 18) {real, imag} */,
  {32'hc1c71048, 32'h41bef18b} /* (5, 22, 17) {real, imag} */,
  {32'hc2a99862, 32'h00000000} /* (5, 22, 16) {real, imag} */,
  {32'hc1c71048, 32'hc1bef18b} /* (5, 22, 15) {real, imag} */,
  {32'h4278778a, 32'h42328223} /* (5, 22, 14) {real, imag} */,
  {32'hbfe0ecb0, 32'hc1c617f6} /* (5, 22, 13) {real, imag} */,
  {32'hc02f04c0, 32'h412f7f18} /* (5, 22, 12) {real, imag} */,
  {32'hc272eea5, 32'hc2084db8} /* (5, 22, 11) {real, imag} */,
  {32'h4232b976, 32'hc23d4d03} /* (5, 22, 10) {real, imag} */,
  {32'hc1d997e7, 32'hc2a36408} /* (5, 22, 9) {real, imag} */,
  {32'hc1ee2d62, 32'h425128e4} /* (5, 22, 8) {real, imag} */,
  {32'h42775e6e, 32'hc103d9a6} /* (5, 22, 7) {real, imag} */,
  {32'h4167edcf, 32'h422c8b1a} /* (5, 22, 6) {real, imag} */,
  {32'h42dc38f9, 32'h429315aa} /* (5, 22, 5) {real, imag} */,
  {32'hc2b581d6, 32'hc2acd972} /* (5, 22, 4) {real, imag} */,
  {32'hc281430e, 32'h433a8b4c} /* (5, 22, 3) {real, imag} */,
  {32'h41832f84, 32'hc2aa38aa} /* (5, 22, 2) {real, imag} */,
  {32'hc3157118, 32'h4371c773} /* (5, 22, 1) {real, imag} */,
  {32'h44585d0a, 32'h00000000} /* (5, 22, 0) {real, imag} */,
  {32'hc3054d6b, 32'hc2eef332} /* (5, 21, 31) {real, imag} */,
  {32'hc2905456, 32'h41c6dc24} /* (5, 21, 30) {real, imag} */,
  {32'h421904b2, 32'hc30d5a76} /* (5, 21, 29) {real, imag} */,
  {32'hc2cdb4a4, 32'h41f7978c} /* (5, 21, 28) {real, imag} */,
  {32'h3f7de6e0, 32'hc1824c1a} /* (5, 21, 27) {real, imag} */,
  {32'hc2f229d4, 32'hc1feabc6} /* (5, 21, 26) {real, imag} */,
  {32'h42c02ea8, 32'h42e3f915} /* (5, 21, 25) {real, imag} */,
  {32'hc2128fd2, 32'hc301d1b3} /* (5, 21, 24) {real, imag} */,
  {32'h3f443880, 32'h421cc1ec} /* (5, 21, 23) {real, imag} */,
  {32'hc0f4c75c, 32'h41efbd7b} /* (5, 21, 22) {real, imag} */,
  {32'hc1003410, 32'hc2b82dcf} /* (5, 21, 21) {real, imag} */,
  {32'h41cd4bee, 32'h410ff798} /* (5, 21, 20) {real, imag} */,
  {32'h3f2b3440, 32'hc1e6d63e} /* (5, 21, 19) {real, imag} */,
  {32'hc1b748b4, 32'h4264f74d} /* (5, 21, 18) {real, imag} */,
  {32'h407eda70, 32'h428fc7f0} /* (5, 21, 17) {real, imag} */,
  {32'h41978d92, 32'h00000000} /* (5, 21, 16) {real, imag} */,
  {32'h407eda70, 32'hc28fc7f0} /* (5, 21, 15) {real, imag} */,
  {32'hc1b748b4, 32'hc264f74d} /* (5, 21, 14) {real, imag} */,
  {32'h3f2b3440, 32'h41e6d63e} /* (5, 21, 13) {real, imag} */,
  {32'h41cd4bee, 32'hc10ff798} /* (5, 21, 12) {real, imag} */,
  {32'hc1003410, 32'h42b82dcf} /* (5, 21, 11) {real, imag} */,
  {32'hc0f4c75c, 32'hc1efbd7b} /* (5, 21, 10) {real, imag} */,
  {32'h3f443880, 32'hc21cc1ec} /* (5, 21, 9) {real, imag} */,
  {32'hc2128fd2, 32'h4301d1b3} /* (5, 21, 8) {real, imag} */,
  {32'h42c02ea8, 32'hc2e3f915} /* (5, 21, 7) {real, imag} */,
  {32'hc2f229d4, 32'h41feabc6} /* (5, 21, 6) {real, imag} */,
  {32'h3f7de6e0, 32'h41824c1a} /* (5, 21, 5) {real, imag} */,
  {32'hc2cdb4a4, 32'hc1f7978c} /* (5, 21, 4) {real, imag} */,
  {32'h421904b2, 32'h430d5a76} /* (5, 21, 3) {real, imag} */,
  {32'hc2905456, 32'hc1c6dc24} /* (5, 21, 2) {real, imag} */,
  {32'hc3054d6b, 32'h42eef332} /* (5, 21, 1) {real, imag} */,
  {32'h44403f92, 32'h00000000} /* (5, 21, 0) {real, imag} */,
  {32'hc25c613c, 32'hc2279a8d} /* (5, 20, 31) {real, imag} */,
  {32'hc2b55a0d, 32'h4122c6c4} /* (5, 20, 30) {real, imag} */,
  {32'h421e9ef8, 32'hc311a847} /* (5, 20, 29) {real, imag} */,
  {32'hc2703a2c, 32'hc2942f89} /* (5, 20, 28) {real, imag} */,
  {32'hc2918444, 32'hc2729eb2} /* (5, 20, 27) {real, imag} */,
  {32'h41c7f7b8, 32'hc1878b18} /* (5, 20, 26) {real, imag} */,
  {32'h41dd9244, 32'h434e3271} /* (5, 20, 25) {real, imag} */,
  {32'hc2d5998e, 32'h41d2825d} /* (5, 20, 24) {real, imag} */,
  {32'hc18ab74c, 32'hc21a317b} /* (5, 20, 23) {real, imag} */,
  {32'hc2de1c92, 32'hc208b17d} /* (5, 20, 22) {real, imag} */,
  {32'hc2339b07, 32'h42c9d7a0} /* (5, 20, 21) {real, imag} */,
  {32'hc1a4e700, 32'hc050f060} /* (5, 20, 20) {real, imag} */,
  {32'h42e99ede, 32'h42167a7d} /* (5, 20, 19) {real, imag} */,
  {32'h4169fcb6, 32'h424e108f} /* (5, 20, 18) {real, imag} */,
  {32'hc20d9d32, 32'hc0594530} /* (5, 20, 17) {real, imag} */,
  {32'hc1e89335, 32'h00000000} /* (5, 20, 16) {real, imag} */,
  {32'hc20d9d32, 32'h40594530} /* (5, 20, 15) {real, imag} */,
  {32'h4169fcb6, 32'hc24e108f} /* (5, 20, 14) {real, imag} */,
  {32'h42e99ede, 32'hc2167a7d} /* (5, 20, 13) {real, imag} */,
  {32'hc1a4e700, 32'h4050f060} /* (5, 20, 12) {real, imag} */,
  {32'hc2339b07, 32'hc2c9d7a0} /* (5, 20, 11) {real, imag} */,
  {32'hc2de1c92, 32'h4208b17d} /* (5, 20, 10) {real, imag} */,
  {32'hc18ab74c, 32'h421a317b} /* (5, 20, 9) {real, imag} */,
  {32'hc2d5998e, 32'hc1d2825d} /* (5, 20, 8) {real, imag} */,
  {32'h41dd9244, 32'hc34e3271} /* (5, 20, 7) {real, imag} */,
  {32'h41c7f7b8, 32'h41878b18} /* (5, 20, 6) {real, imag} */,
  {32'hc2918444, 32'h42729eb2} /* (5, 20, 5) {real, imag} */,
  {32'hc2703a2c, 32'h42942f89} /* (5, 20, 4) {real, imag} */,
  {32'h421e9ef8, 32'h4311a847} /* (5, 20, 3) {real, imag} */,
  {32'hc2b55a0d, 32'hc122c6c4} /* (5, 20, 2) {real, imag} */,
  {32'hc25c613c, 32'h42279a8d} /* (5, 20, 1) {real, imag} */,
  {32'h444612eb, 32'h00000000} /* (5, 20, 0) {real, imag} */,
  {32'hc33a1410, 32'hc1ab89a8} /* (5, 19, 31) {real, imag} */,
  {32'hc2aa292e, 32'hc236ed44} /* (5, 19, 30) {real, imag} */,
  {32'hc1978d00, 32'hc31d8f8a} /* (5, 19, 29) {real, imag} */,
  {32'hc2b0cf86, 32'hc275a038} /* (5, 19, 28) {real, imag} */,
  {32'hc276ce49, 32'hc2511d7a} /* (5, 19, 27) {real, imag} */,
  {32'h41ec5304, 32'h420120a3} /* (5, 19, 26) {real, imag} */,
  {32'h42e45732, 32'h41cacf12} /* (5, 19, 25) {real, imag} */,
  {32'hc2d11fd0, 32'h41b4fee0} /* (5, 19, 24) {real, imag} */,
  {32'hc2c0c84c, 32'hc1800e70} /* (5, 19, 23) {real, imag} */,
  {32'hc22cbd86, 32'hbef8b800} /* (5, 19, 22) {real, imag} */,
  {32'hc2c7d986, 32'h426c02aa} /* (5, 19, 21) {real, imag} */,
  {32'hc2bce2bd, 32'h412ea6e8} /* (5, 19, 20) {real, imag} */,
  {32'hc22b8fa9, 32'hc1d3ee7c} /* (5, 19, 19) {real, imag} */,
  {32'hbfc725c0, 32'h419c2184} /* (5, 19, 18) {real, imag} */,
  {32'h4190534a, 32'h422792dc} /* (5, 19, 17) {real, imag} */,
  {32'h4067d948, 32'h00000000} /* (5, 19, 16) {real, imag} */,
  {32'h4190534a, 32'hc22792dc} /* (5, 19, 15) {real, imag} */,
  {32'hbfc725c0, 32'hc19c2184} /* (5, 19, 14) {real, imag} */,
  {32'hc22b8fa9, 32'h41d3ee7c} /* (5, 19, 13) {real, imag} */,
  {32'hc2bce2bd, 32'hc12ea6e8} /* (5, 19, 12) {real, imag} */,
  {32'hc2c7d986, 32'hc26c02aa} /* (5, 19, 11) {real, imag} */,
  {32'hc22cbd86, 32'h3ef8b800} /* (5, 19, 10) {real, imag} */,
  {32'hc2c0c84c, 32'h41800e70} /* (5, 19, 9) {real, imag} */,
  {32'hc2d11fd0, 32'hc1b4fee0} /* (5, 19, 8) {real, imag} */,
  {32'h42e45732, 32'hc1cacf12} /* (5, 19, 7) {real, imag} */,
  {32'h41ec5304, 32'hc20120a3} /* (5, 19, 6) {real, imag} */,
  {32'hc276ce49, 32'h42511d7a} /* (5, 19, 5) {real, imag} */,
  {32'hc2b0cf86, 32'h4275a038} /* (5, 19, 4) {real, imag} */,
  {32'hc1978d00, 32'h431d8f8a} /* (5, 19, 3) {real, imag} */,
  {32'hc2aa292e, 32'h4236ed44} /* (5, 19, 2) {real, imag} */,
  {32'hc33a1410, 32'h41ab89a8} /* (5, 19, 1) {real, imag} */,
  {32'h43921b0c, 32'h00000000} /* (5, 19, 0) {real, imag} */,
  {32'hc3871ec2, 32'h41ad5516} /* (5, 18, 31) {real, imag} */,
  {32'hc1cb931c, 32'h42c65f19} /* (5, 18, 30) {real, imag} */,
  {32'hc285b697, 32'hc306b288} /* (5, 18, 29) {real, imag} */,
  {32'hc3093d40, 32'hc2b7884b} /* (5, 18, 28) {real, imag} */,
  {32'h4288f802, 32'hc155ef58} /* (5, 18, 27) {real, imag} */,
  {32'h41816de6, 32'h418f2306} /* (5, 18, 26) {real, imag} */,
  {32'h422e85f4, 32'h41b133e4} /* (5, 18, 25) {real, imag} */,
  {32'h406002c0, 32'h428bc79d} /* (5, 18, 24) {real, imag} */,
  {32'h424e0adc, 32'h4280f9ce} /* (5, 18, 23) {real, imag} */,
  {32'h407734ec, 32'hc080dfd0} /* (5, 18, 22) {real, imag} */,
  {32'h42008844, 32'hc17db6fc} /* (5, 18, 21) {real, imag} */,
  {32'hc2dc6b40, 32'hc1c439fd} /* (5, 18, 20) {real, imag} */,
  {32'hc1cdaf28, 32'h42942408} /* (5, 18, 19) {real, imag} */,
  {32'hc30bceed, 32'h41affbfa} /* (5, 18, 18) {real, imag} */,
  {32'hc1eb9f3a, 32'h4289febc} /* (5, 18, 17) {real, imag} */,
  {32'hc2ac5c58, 32'h00000000} /* (5, 18, 16) {real, imag} */,
  {32'hc1eb9f3a, 32'hc289febc} /* (5, 18, 15) {real, imag} */,
  {32'hc30bceed, 32'hc1affbfa} /* (5, 18, 14) {real, imag} */,
  {32'hc1cdaf28, 32'hc2942408} /* (5, 18, 13) {real, imag} */,
  {32'hc2dc6b40, 32'h41c439fd} /* (5, 18, 12) {real, imag} */,
  {32'h42008844, 32'h417db6fc} /* (5, 18, 11) {real, imag} */,
  {32'h407734ec, 32'h4080dfd0} /* (5, 18, 10) {real, imag} */,
  {32'h424e0adc, 32'hc280f9ce} /* (5, 18, 9) {real, imag} */,
  {32'h406002c0, 32'hc28bc79d} /* (5, 18, 8) {real, imag} */,
  {32'h422e85f4, 32'hc1b133e4} /* (5, 18, 7) {real, imag} */,
  {32'h41816de6, 32'hc18f2306} /* (5, 18, 6) {real, imag} */,
  {32'h4288f802, 32'h4155ef58} /* (5, 18, 5) {real, imag} */,
  {32'hc3093d40, 32'h42b7884b} /* (5, 18, 4) {real, imag} */,
  {32'hc285b697, 32'h4306b288} /* (5, 18, 3) {real, imag} */,
  {32'hc1cb931c, 32'hc2c65f19} /* (5, 18, 2) {real, imag} */,
  {32'hc3871ec2, 32'hc1ad5516} /* (5, 18, 1) {real, imag} */,
  {32'h42131c80, 32'h00000000} /* (5, 18, 0) {real, imag} */,
  {32'hc3d87e0f, 32'h40d755a0} /* (5, 17, 31) {real, imag} */,
  {32'h41d7f229, 32'h430e05ea} /* (5, 17, 30) {real, imag} */,
  {32'h41d00589, 32'h422c034e} /* (5, 17, 29) {real, imag} */,
  {32'h42600416, 32'hc10c7da4} /* (5, 17, 28) {real, imag} */,
  {32'h418a2c08, 32'h42ae17ac} /* (5, 17, 27) {real, imag} */,
  {32'h405d54e0, 32'hc2b2a34b} /* (5, 17, 26) {real, imag} */,
  {32'hc282f3d4, 32'h4214c586} /* (5, 17, 25) {real, imag} */,
  {32'h40d31f3c, 32'h41fd69fc} /* (5, 17, 24) {real, imag} */,
  {32'hc23a368f, 32'h4207f064} /* (5, 17, 23) {real, imag} */,
  {32'h41abe4cc, 32'h41b1a918} /* (5, 17, 22) {real, imag} */,
  {32'hc210cbde, 32'hc13a43c8} /* (5, 17, 21) {real, imag} */,
  {32'h41b13e88, 32'h4220feee} /* (5, 17, 20) {real, imag} */,
  {32'h40b47600, 32'h423c0ae1} /* (5, 17, 19) {real, imag} */,
  {32'h41626b1f, 32'hc0d679a8} /* (5, 17, 18) {real, imag} */,
  {32'hc25f17b9, 32'hc1ff65fd} /* (5, 17, 17) {real, imag} */,
  {32'h426f0d12, 32'h00000000} /* (5, 17, 16) {real, imag} */,
  {32'hc25f17b9, 32'h41ff65fd} /* (5, 17, 15) {real, imag} */,
  {32'h41626b1f, 32'h40d679a8} /* (5, 17, 14) {real, imag} */,
  {32'h40b47600, 32'hc23c0ae1} /* (5, 17, 13) {real, imag} */,
  {32'h41b13e88, 32'hc220feee} /* (5, 17, 12) {real, imag} */,
  {32'hc210cbde, 32'h413a43c8} /* (5, 17, 11) {real, imag} */,
  {32'h41abe4cc, 32'hc1b1a918} /* (5, 17, 10) {real, imag} */,
  {32'hc23a368f, 32'hc207f064} /* (5, 17, 9) {real, imag} */,
  {32'h40d31f3c, 32'hc1fd69fc} /* (5, 17, 8) {real, imag} */,
  {32'hc282f3d4, 32'hc214c586} /* (5, 17, 7) {real, imag} */,
  {32'h405d54e0, 32'h42b2a34b} /* (5, 17, 6) {real, imag} */,
  {32'h418a2c08, 32'hc2ae17ac} /* (5, 17, 5) {real, imag} */,
  {32'h42600416, 32'h410c7da4} /* (5, 17, 4) {real, imag} */,
  {32'h41d00589, 32'hc22c034e} /* (5, 17, 3) {real, imag} */,
  {32'h41d7f229, 32'hc30e05ea} /* (5, 17, 2) {real, imag} */,
  {32'hc3d87e0f, 32'hc0d755a0} /* (5, 17, 1) {real, imag} */,
  {32'hc2851e74, 32'h00000000} /* (5, 17, 0) {real, imag} */,
  {32'hc3f9e8eb, 32'hc2cc97d6} /* (5, 16, 31) {real, imag} */,
  {32'hc2c35311, 32'h42caddd0} /* (5, 16, 30) {real, imag} */,
  {32'h427ef099, 32'hc1b1479c} /* (5, 16, 29) {real, imag} */,
  {32'h40f916c8, 32'hc2c0cd62} /* (5, 16, 28) {real, imag} */,
  {32'h42e3eee3, 32'h4220a392} /* (5, 16, 27) {real, imag} */,
  {32'hc1f62a0a, 32'hbfaf1058} /* (5, 16, 26) {real, imag} */,
  {32'h432eec83, 32'hc12ac17e} /* (5, 16, 25) {real, imag} */,
  {32'hc22210d8, 32'h424811f0} /* (5, 16, 24) {real, imag} */,
  {32'h42683723, 32'hc226b36a} /* (5, 16, 23) {real, imag} */,
  {32'hc20030c5, 32'h42a54472} /* (5, 16, 22) {real, imag} */,
  {32'hc258cfad, 32'hc2a0bf86} /* (5, 16, 21) {real, imag} */,
  {32'hc2811e3e, 32'hc13324af} /* (5, 16, 20) {real, imag} */,
  {32'h41521868, 32'h424fb3cb} /* (5, 16, 19) {real, imag} */,
  {32'hc13ca89a, 32'h414b9364} /* (5, 16, 18) {real, imag} */,
  {32'h426301e1, 32'hc2286e2a} /* (5, 16, 17) {real, imag} */,
  {32'hc09111bc, 32'h00000000} /* (5, 16, 16) {real, imag} */,
  {32'h426301e1, 32'h42286e2a} /* (5, 16, 15) {real, imag} */,
  {32'hc13ca89a, 32'hc14b9364} /* (5, 16, 14) {real, imag} */,
  {32'h41521868, 32'hc24fb3cb} /* (5, 16, 13) {real, imag} */,
  {32'hc2811e3e, 32'h413324af} /* (5, 16, 12) {real, imag} */,
  {32'hc258cfad, 32'h42a0bf86} /* (5, 16, 11) {real, imag} */,
  {32'hc20030c5, 32'hc2a54472} /* (5, 16, 10) {real, imag} */,
  {32'h42683723, 32'h4226b36a} /* (5, 16, 9) {real, imag} */,
  {32'hc22210d8, 32'hc24811f0} /* (5, 16, 8) {real, imag} */,
  {32'h432eec83, 32'h412ac17e} /* (5, 16, 7) {real, imag} */,
  {32'hc1f62a0a, 32'h3faf1058} /* (5, 16, 6) {real, imag} */,
  {32'h42e3eee3, 32'hc220a392} /* (5, 16, 5) {real, imag} */,
  {32'h40f916c8, 32'h42c0cd62} /* (5, 16, 4) {real, imag} */,
  {32'h427ef099, 32'h41b1479c} /* (5, 16, 3) {real, imag} */,
  {32'hc2c35311, 32'hc2caddd0} /* (5, 16, 2) {real, imag} */,
  {32'hc3f9e8eb, 32'h42cc97d6} /* (5, 16, 1) {real, imag} */,
  {32'hc30e7064, 32'h00000000} /* (5, 16, 0) {real, imag} */,
  {32'hc3ceea47, 32'hc36888ef} /* (5, 15, 31) {real, imag} */,
  {32'h402b42f8, 32'h42e7da21} /* (5, 15, 30) {real, imag} */,
  {32'h423f6adc, 32'hc3693328} /* (5, 15, 29) {real, imag} */,
  {32'h428d4ec9, 32'hc1a6e0e2} /* (5, 15, 28) {real, imag} */,
  {32'hc1ac2662, 32'h416a07b0} /* (5, 15, 27) {real, imag} */,
  {32'h42a0ae6b, 32'hc20e6d96} /* (5, 15, 26) {real, imag} */,
  {32'h42b5019c, 32'h4271c8a2} /* (5, 15, 25) {real, imag} */,
  {32'h3fb47970, 32'h40849c78} /* (5, 15, 24) {real, imag} */,
  {32'hc29f2f7a, 32'h4112412a} /* (5, 15, 23) {real, imag} */,
  {32'hc1178899, 32'h429eb7cb} /* (5, 15, 22) {real, imag} */,
  {32'h42251f94, 32'hc282afd5} /* (5, 15, 21) {real, imag} */,
  {32'hc20d9d71, 32'h42b22f71} /* (5, 15, 20) {real, imag} */,
  {32'hc3113a63, 32'hc296c4af} /* (5, 15, 19) {real, imag} */,
  {32'h410688ab, 32'hc1b7c78e} /* (5, 15, 18) {real, imag} */,
  {32'hc2abbb44, 32'h42666d12} /* (5, 15, 17) {real, imag} */,
  {32'hc227d99e, 32'h00000000} /* (5, 15, 16) {real, imag} */,
  {32'hc2abbb44, 32'hc2666d12} /* (5, 15, 15) {real, imag} */,
  {32'h410688ab, 32'h41b7c78e} /* (5, 15, 14) {real, imag} */,
  {32'hc3113a63, 32'h4296c4af} /* (5, 15, 13) {real, imag} */,
  {32'hc20d9d71, 32'hc2b22f71} /* (5, 15, 12) {real, imag} */,
  {32'h42251f94, 32'h4282afd5} /* (5, 15, 11) {real, imag} */,
  {32'hc1178899, 32'hc29eb7cb} /* (5, 15, 10) {real, imag} */,
  {32'hc29f2f7a, 32'hc112412a} /* (5, 15, 9) {real, imag} */,
  {32'h3fb47970, 32'hc0849c78} /* (5, 15, 8) {real, imag} */,
  {32'h42b5019c, 32'hc271c8a2} /* (5, 15, 7) {real, imag} */,
  {32'h42a0ae6b, 32'h420e6d96} /* (5, 15, 6) {real, imag} */,
  {32'hc1ac2662, 32'hc16a07b0} /* (5, 15, 5) {real, imag} */,
  {32'h428d4ec9, 32'h41a6e0e2} /* (5, 15, 4) {real, imag} */,
  {32'h423f6adc, 32'h43693328} /* (5, 15, 3) {real, imag} */,
  {32'h402b42f8, 32'hc2e7da21} /* (5, 15, 2) {real, imag} */,
  {32'hc3ceea47, 32'h436888ef} /* (5, 15, 1) {real, imag} */,
  {32'hc3e65a8f, 32'h00000000} /* (5, 15, 0) {real, imag} */,
  {32'hc3a66182, 32'hc2bd5c0e} /* (5, 14, 31) {real, imag} */,
  {32'h4227657e, 32'hc2f14d77} /* (5, 14, 30) {real, imag} */,
  {32'h42a8986d, 32'hc31b2330} /* (5, 14, 29) {real, imag} */,
  {32'h41513438, 32'hc2df6273} /* (5, 14, 28) {real, imag} */,
  {32'hc23c8f1a, 32'h4292f208} /* (5, 14, 27) {real, imag} */,
  {32'h4234e47c, 32'hc007a950} /* (5, 14, 26) {real, imag} */,
  {32'h4261e8cc, 32'hc271141a} /* (5, 14, 25) {real, imag} */,
  {32'hc0817610, 32'hc2874403} /* (5, 14, 24) {real, imag} */,
  {32'h3fbc9e40, 32'h42cbbaf2} /* (5, 14, 23) {real, imag} */,
  {32'hc09c63b6, 32'hc2887c4d} /* (5, 14, 22) {real, imag} */,
  {32'h42b5ed72, 32'h429b05dc} /* (5, 14, 21) {real, imag} */,
  {32'h42312329, 32'h41029a16} /* (5, 14, 20) {real, imag} */,
  {32'hc229543e, 32'h4177dfd4} /* (5, 14, 19) {real, imag} */,
  {32'h429c9ab8, 32'h401468e0} /* (5, 14, 18) {real, imag} */,
  {32'hc276454b, 32'hc20f5ba3} /* (5, 14, 17) {real, imag} */,
  {32'h428684cc, 32'h00000000} /* (5, 14, 16) {real, imag} */,
  {32'hc276454b, 32'h420f5ba3} /* (5, 14, 15) {real, imag} */,
  {32'h429c9ab8, 32'hc01468e0} /* (5, 14, 14) {real, imag} */,
  {32'hc229543e, 32'hc177dfd4} /* (5, 14, 13) {real, imag} */,
  {32'h42312329, 32'hc1029a16} /* (5, 14, 12) {real, imag} */,
  {32'h42b5ed72, 32'hc29b05dc} /* (5, 14, 11) {real, imag} */,
  {32'hc09c63b6, 32'h42887c4d} /* (5, 14, 10) {real, imag} */,
  {32'h3fbc9e40, 32'hc2cbbaf2} /* (5, 14, 9) {real, imag} */,
  {32'hc0817610, 32'h42874403} /* (5, 14, 8) {real, imag} */,
  {32'h4261e8cc, 32'h4271141a} /* (5, 14, 7) {real, imag} */,
  {32'h4234e47c, 32'h4007a950} /* (5, 14, 6) {real, imag} */,
  {32'hc23c8f1a, 32'hc292f208} /* (5, 14, 5) {real, imag} */,
  {32'h41513438, 32'h42df6273} /* (5, 14, 4) {real, imag} */,
  {32'h42a8986d, 32'h431b2330} /* (5, 14, 3) {real, imag} */,
  {32'h4227657e, 32'h42f14d77} /* (5, 14, 2) {real, imag} */,
  {32'hc3a66182, 32'h42bd5c0e} /* (5, 14, 1) {real, imag} */,
  {32'hc421ceac, 32'h00000000} /* (5, 14, 0) {real, imag} */,
  {32'hc2901a60, 32'hc35fbf49} /* (5, 13, 31) {real, imag} */,
  {32'hc1a0dd72, 32'hc36c444d} /* (5, 13, 30) {real, imag} */,
  {32'h42cf1bd8, 32'hc2232b3a} /* (5, 13, 29) {real, imag} */,
  {32'hc2933a6a, 32'hc31f59ee} /* (5, 13, 28) {real, imag} */,
  {32'hc2b51ca2, 32'h43475f9e} /* (5, 13, 27) {real, imag} */,
  {32'h43454778, 32'h42e56574} /* (5, 13, 26) {real, imag} */,
  {32'h42608ecf, 32'hc25435dd} /* (5, 13, 25) {real, imag} */,
  {32'hc2a7f81e, 32'h418ca934} /* (5, 13, 24) {real, imag} */,
  {32'h42642a71, 32'h42a6ff7e} /* (5, 13, 23) {real, imag} */,
  {32'h41b16f6c, 32'hc2e3da4c} /* (5, 13, 22) {real, imag} */,
  {32'hc2968342, 32'h3f74c8a0} /* (5, 13, 21) {real, imag} */,
  {32'h423f306e, 32'hc0ebe530} /* (5, 13, 20) {real, imag} */,
  {32'hc287c768, 32'hc2c6f4bf} /* (5, 13, 19) {real, imag} */,
  {32'hc23cfc24, 32'h4283325e} /* (5, 13, 18) {real, imag} */,
  {32'h425556ef, 32'hc20b89fa} /* (5, 13, 17) {real, imag} */,
  {32'hc1573bd6, 32'h00000000} /* (5, 13, 16) {real, imag} */,
  {32'h425556ef, 32'h420b89fa} /* (5, 13, 15) {real, imag} */,
  {32'hc23cfc24, 32'hc283325e} /* (5, 13, 14) {real, imag} */,
  {32'hc287c768, 32'h42c6f4bf} /* (5, 13, 13) {real, imag} */,
  {32'h423f306e, 32'h40ebe530} /* (5, 13, 12) {real, imag} */,
  {32'hc2968342, 32'hbf74c8a0} /* (5, 13, 11) {real, imag} */,
  {32'h41b16f6c, 32'h42e3da4c} /* (5, 13, 10) {real, imag} */,
  {32'h42642a71, 32'hc2a6ff7e} /* (5, 13, 9) {real, imag} */,
  {32'hc2a7f81e, 32'hc18ca934} /* (5, 13, 8) {real, imag} */,
  {32'h42608ecf, 32'h425435dd} /* (5, 13, 7) {real, imag} */,
  {32'h43454778, 32'hc2e56574} /* (5, 13, 6) {real, imag} */,
  {32'hc2b51ca2, 32'hc3475f9e} /* (5, 13, 5) {real, imag} */,
  {32'hc2933a6a, 32'h431f59ee} /* (5, 13, 4) {real, imag} */,
  {32'h42cf1bd8, 32'h42232b3a} /* (5, 13, 3) {real, imag} */,
  {32'hc1a0dd72, 32'h436c444d} /* (5, 13, 2) {real, imag} */,
  {32'hc2901a60, 32'h435fbf49} /* (5, 13, 1) {real, imag} */,
  {32'hc3f17ebc, 32'h00000000} /* (5, 13, 0) {real, imag} */,
  {32'h42881c4e, 32'hc2f32dae} /* (5, 12, 31) {real, imag} */,
  {32'h431065e0, 32'hc305f511} /* (5, 12, 30) {real, imag} */,
  {32'h430aa958, 32'h4286d878} /* (5, 12, 29) {real, imag} */,
  {32'hc29b5092, 32'hc20c787e} /* (5, 12, 28) {real, imag} */,
  {32'hc3031fa4, 32'h42f1c2df} /* (5, 12, 27) {real, imag} */,
  {32'h42efbd0e, 32'h430b108d} /* (5, 12, 26) {real, imag} */,
  {32'hc2ab9f7b, 32'hc11f0d40} /* (5, 12, 25) {real, imag} */,
  {32'h423902d7, 32'h4289cc2d} /* (5, 12, 24) {real, imag} */,
  {32'h4239087b, 32'hc0832910} /* (5, 12, 23) {real, imag} */,
  {32'hc24e4b25, 32'hc27894bf} /* (5, 12, 22) {real, imag} */,
  {32'hc155b2c4, 32'h3f1b7700} /* (5, 12, 21) {real, imag} */,
  {32'hc1b730d8, 32'hc2b77e05} /* (5, 12, 20) {real, imag} */,
  {32'h41ab4548, 32'h4298a5d8} /* (5, 12, 19) {real, imag} */,
  {32'h3e727280, 32'hc1e2ef62} /* (5, 12, 18) {real, imag} */,
  {32'hc10f014e, 32'hc29572ba} /* (5, 12, 17) {real, imag} */,
  {32'hc2b11d75, 32'h00000000} /* (5, 12, 16) {real, imag} */,
  {32'hc10f014e, 32'h429572ba} /* (5, 12, 15) {real, imag} */,
  {32'h3e727280, 32'h41e2ef62} /* (5, 12, 14) {real, imag} */,
  {32'h41ab4548, 32'hc298a5d8} /* (5, 12, 13) {real, imag} */,
  {32'hc1b730d8, 32'h42b77e05} /* (5, 12, 12) {real, imag} */,
  {32'hc155b2c4, 32'hbf1b7700} /* (5, 12, 11) {real, imag} */,
  {32'hc24e4b25, 32'h427894bf} /* (5, 12, 10) {real, imag} */,
  {32'h4239087b, 32'h40832910} /* (5, 12, 9) {real, imag} */,
  {32'h423902d7, 32'hc289cc2d} /* (5, 12, 8) {real, imag} */,
  {32'hc2ab9f7b, 32'h411f0d40} /* (5, 12, 7) {real, imag} */,
  {32'h42efbd0e, 32'hc30b108d} /* (5, 12, 6) {real, imag} */,
  {32'hc3031fa4, 32'hc2f1c2df} /* (5, 12, 5) {real, imag} */,
  {32'hc29b5092, 32'h420c787e} /* (5, 12, 4) {real, imag} */,
  {32'h430aa958, 32'hc286d878} /* (5, 12, 3) {real, imag} */,
  {32'h431065e0, 32'h4305f511} /* (5, 12, 2) {real, imag} */,
  {32'h42881c4e, 32'h42f32dae} /* (5, 12, 1) {real, imag} */,
  {32'hc3123ac4, 32'h00000000} /* (5, 12, 0) {real, imag} */,
  {32'h431e4923, 32'hc39c77f6} /* (5, 11, 31) {real, imag} */,
  {32'h42996248, 32'hc25b77be} /* (5, 11, 30) {real, imag} */,
  {32'h4349dc36, 32'h420599f6} /* (5, 11, 29) {real, imag} */,
  {32'h4266896b, 32'hc284e717} /* (5, 11, 28) {real, imag} */,
  {32'hc206f428, 32'h42cd19ac} /* (5, 11, 27) {real, imag} */,
  {32'h431c1a94, 32'h40d91450} /* (5, 11, 26) {real, imag} */,
  {32'hc0ba8b98, 32'h4210dc32} /* (5, 11, 25) {real, imag} */,
  {32'h4142ce88, 32'h4237888c} /* (5, 11, 24) {real, imag} */,
  {32'h4304636e, 32'h42b0f99a} /* (5, 11, 23) {real, imag} */,
  {32'hc2664bba, 32'h423677e2} /* (5, 11, 22) {real, imag} */,
  {32'hc2b3b7e0, 32'h42aeffb1} /* (5, 11, 21) {real, imag} */,
  {32'hc300a5a5, 32'h42a3e6d5} /* (5, 11, 20) {real, imag} */,
  {32'h420c3067, 32'h426af91f} /* (5, 11, 19) {real, imag} */,
  {32'h426eef92, 32'hc194815e} /* (5, 11, 18) {real, imag} */,
  {32'hc2b3a710, 32'h4222d4de} /* (5, 11, 17) {real, imag} */,
  {32'h42c901f6, 32'h00000000} /* (5, 11, 16) {real, imag} */,
  {32'hc2b3a710, 32'hc222d4de} /* (5, 11, 15) {real, imag} */,
  {32'h426eef92, 32'h4194815e} /* (5, 11, 14) {real, imag} */,
  {32'h420c3067, 32'hc26af91f} /* (5, 11, 13) {real, imag} */,
  {32'hc300a5a5, 32'hc2a3e6d5} /* (5, 11, 12) {real, imag} */,
  {32'hc2b3b7e0, 32'hc2aeffb1} /* (5, 11, 11) {real, imag} */,
  {32'hc2664bba, 32'hc23677e2} /* (5, 11, 10) {real, imag} */,
  {32'h4304636e, 32'hc2b0f99a} /* (5, 11, 9) {real, imag} */,
  {32'h4142ce88, 32'hc237888c} /* (5, 11, 8) {real, imag} */,
  {32'hc0ba8b98, 32'hc210dc32} /* (5, 11, 7) {real, imag} */,
  {32'h431c1a94, 32'hc0d91450} /* (5, 11, 6) {real, imag} */,
  {32'hc206f428, 32'hc2cd19ac} /* (5, 11, 5) {real, imag} */,
  {32'h4266896b, 32'h4284e717} /* (5, 11, 4) {real, imag} */,
  {32'h4349dc36, 32'hc20599f6} /* (5, 11, 3) {real, imag} */,
  {32'h42996248, 32'h425b77be} /* (5, 11, 2) {real, imag} */,
  {32'h431e4923, 32'h439c77f6} /* (5, 11, 1) {real, imag} */,
  {32'h4346d0ba, 32'h00000000} /* (5, 11, 0) {real, imag} */,
  {32'h42cc1dd5, 32'hc3bec316} /* (5, 10, 31) {real, imag} */,
  {32'h42e91543, 32'hc2281a5c} /* (5, 10, 30) {real, imag} */,
  {32'h4296e0c6, 32'hc19c2220} /* (5, 10, 29) {real, imag} */,
  {32'h42433f74, 32'hc2bc8f7a} /* (5, 10, 28) {real, imag} */,
  {32'hc19c3374, 32'h40a38f78} /* (5, 10, 27) {real, imag} */,
  {32'hc230ca1b, 32'hc16f7cd0} /* (5, 10, 26) {real, imag} */,
  {32'h411348c6, 32'hc1323106} /* (5, 10, 25) {real, imag} */,
  {32'h41b7748e, 32'hc36bdb65} /* (5, 10, 24) {real, imag} */,
  {32'hc26b5da0, 32'h434d1d0a} /* (5, 10, 23) {real, imag} */,
  {32'h4297edf5, 32'h42ffbe9e} /* (5, 10, 22) {real, imag} */,
  {32'hc21b9e13, 32'hc2f5f6d4} /* (5, 10, 21) {real, imag} */,
  {32'h42ac785e, 32'h426f292a} /* (5, 10, 20) {real, imag} */,
  {32'h4254f9d8, 32'h41a8b8da} /* (5, 10, 19) {real, imag} */,
  {32'hc216eaec, 32'h42854518} /* (5, 10, 18) {real, imag} */,
  {32'hc107432f, 32'h42349178} /* (5, 10, 17) {real, imag} */,
  {32'hc27682f4, 32'h00000000} /* (5, 10, 16) {real, imag} */,
  {32'hc107432f, 32'hc2349178} /* (5, 10, 15) {real, imag} */,
  {32'hc216eaec, 32'hc2854518} /* (5, 10, 14) {real, imag} */,
  {32'h4254f9d8, 32'hc1a8b8da} /* (5, 10, 13) {real, imag} */,
  {32'h42ac785e, 32'hc26f292a} /* (5, 10, 12) {real, imag} */,
  {32'hc21b9e13, 32'h42f5f6d4} /* (5, 10, 11) {real, imag} */,
  {32'h4297edf5, 32'hc2ffbe9e} /* (5, 10, 10) {real, imag} */,
  {32'hc26b5da0, 32'hc34d1d0a} /* (5, 10, 9) {real, imag} */,
  {32'h41b7748e, 32'h436bdb65} /* (5, 10, 8) {real, imag} */,
  {32'h411348c6, 32'h41323106} /* (5, 10, 7) {real, imag} */,
  {32'hc230ca1b, 32'h416f7cd0} /* (5, 10, 6) {real, imag} */,
  {32'hc19c3374, 32'hc0a38f78} /* (5, 10, 5) {real, imag} */,
  {32'h42433f74, 32'h42bc8f7a} /* (5, 10, 4) {real, imag} */,
  {32'h4296e0c6, 32'h419c2220} /* (5, 10, 3) {real, imag} */,
  {32'h42e91543, 32'h42281a5c} /* (5, 10, 2) {real, imag} */,
  {32'h42cc1dd5, 32'h43bec316} /* (5, 10, 1) {real, imag} */,
  {32'h43a5b66c, 32'h00000000} /* (5, 10, 0) {real, imag} */,
  {32'h429e4805, 32'hc3a6c253} /* (5, 9, 31) {real, imag} */,
  {32'h42be638d, 32'h421b2260} /* (5, 9, 30) {real, imag} */,
  {32'h4279f48e, 32'h41afd17e} /* (5, 9, 29) {real, imag} */,
  {32'h4238a1ec, 32'hc1953085} /* (5, 9, 28) {real, imag} */,
  {32'hc1f382d9, 32'hc20c950d} /* (5, 9, 27) {real, imag} */,
  {32'h4302140a, 32'h423ed4e4} /* (5, 9, 26) {real, imag} */,
  {32'hc223472e, 32'h41f1555a} /* (5, 9, 25) {real, imag} */,
  {32'h42332f1a, 32'hc2a7078a} /* (5, 9, 24) {real, imag} */,
  {32'h410de37a, 32'h4286fa36} /* (5, 9, 23) {real, imag} */,
  {32'h42e71e5d, 32'hc1a19a8b} /* (5, 9, 22) {real, imag} */,
  {32'h41d57e22, 32'h40c18110} /* (5, 9, 21) {real, imag} */,
  {32'hc2c18fc9, 32'hc1e96618} /* (5, 9, 20) {real, imag} */,
  {32'hc254d48d, 32'h42697bdc} /* (5, 9, 19) {real, imag} */,
  {32'h423c0333, 32'hc25f5362} /* (5, 9, 18) {real, imag} */,
  {32'h420b3909, 32'h42577b66} /* (5, 9, 17) {real, imag} */,
  {32'hc2a3cc98, 32'h00000000} /* (5, 9, 16) {real, imag} */,
  {32'h420b3909, 32'hc2577b66} /* (5, 9, 15) {real, imag} */,
  {32'h423c0333, 32'h425f5362} /* (5, 9, 14) {real, imag} */,
  {32'hc254d48d, 32'hc2697bdc} /* (5, 9, 13) {real, imag} */,
  {32'hc2c18fc9, 32'h41e96618} /* (5, 9, 12) {real, imag} */,
  {32'h41d57e22, 32'hc0c18110} /* (5, 9, 11) {real, imag} */,
  {32'h42e71e5d, 32'h41a19a8b} /* (5, 9, 10) {real, imag} */,
  {32'h410de37a, 32'hc286fa36} /* (5, 9, 9) {real, imag} */,
  {32'h42332f1a, 32'h42a7078a} /* (5, 9, 8) {real, imag} */,
  {32'hc223472e, 32'hc1f1555a} /* (5, 9, 7) {real, imag} */,
  {32'h4302140a, 32'hc23ed4e4} /* (5, 9, 6) {real, imag} */,
  {32'hc1f382d9, 32'h420c950d} /* (5, 9, 5) {real, imag} */,
  {32'h4238a1ec, 32'h41953085} /* (5, 9, 4) {real, imag} */,
  {32'h4279f48e, 32'hc1afd17e} /* (5, 9, 3) {real, imag} */,
  {32'h42be638d, 32'hc21b2260} /* (5, 9, 2) {real, imag} */,
  {32'h429e4805, 32'h43a6c253} /* (5, 9, 1) {real, imag} */,
  {32'h442c0ed7, 32'h00000000} /* (5, 9, 0) {real, imag} */,
  {32'h43281039, 32'hc3ccec91} /* (5, 8, 31) {real, imag} */,
  {32'h431e2e54, 32'h4393dd65} /* (5, 8, 30) {real, imag} */,
  {32'h43598d04, 32'hc2d0d8be} /* (5, 8, 29) {real, imag} */,
  {32'h428f4622, 32'h426ef0dc} /* (5, 8, 28) {real, imag} */,
  {32'hc297f78d, 32'hc16f8574} /* (5, 8, 27) {real, imag} */,
  {32'h42323977, 32'h4215c822} /* (5, 8, 26) {real, imag} */,
  {32'hc2360250, 32'h426f3d3e} /* (5, 8, 25) {real, imag} */,
  {32'h41a9e1ba, 32'hc30f8c8f} /* (5, 8, 24) {real, imag} */,
  {32'h420e2ab9, 32'h41958d5c} /* (5, 8, 23) {real, imag} */,
  {32'hc2c11280, 32'h42b43374} /* (5, 8, 22) {real, imag} */,
  {32'h42da8d51, 32'h40aee4bc} /* (5, 8, 21) {real, imag} */,
  {32'h41b52bf0, 32'hc246b73c} /* (5, 8, 20) {real, imag} */,
  {32'hc2260b85, 32'hc205b1f8} /* (5, 8, 19) {real, imag} */,
  {32'hc29d990a, 32'hc02925d0} /* (5, 8, 18) {real, imag} */,
  {32'hc1693063, 32'hc16667f6} /* (5, 8, 17) {real, imag} */,
  {32'hc28d6063, 32'h00000000} /* (5, 8, 16) {real, imag} */,
  {32'hc1693063, 32'h416667f6} /* (5, 8, 15) {real, imag} */,
  {32'hc29d990a, 32'h402925d0} /* (5, 8, 14) {real, imag} */,
  {32'hc2260b85, 32'h4205b1f8} /* (5, 8, 13) {real, imag} */,
  {32'h41b52bf0, 32'h4246b73c} /* (5, 8, 12) {real, imag} */,
  {32'h42da8d51, 32'hc0aee4bc} /* (5, 8, 11) {real, imag} */,
  {32'hc2c11280, 32'hc2b43374} /* (5, 8, 10) {real, imag} */,
  {32'h420e2ab9, 32'hc1958d5c} /* (5, 8, 9) {real, imag} */,
  {32'h41a9e1ba, 32'h430f8c8f} /* (5, 8, 8) {real, imag} */,
  {32'hc2360250, 32'hc26f3d3e} /* (5, 8, 7) {real, imag} */,
  {32'h42323977, 32'hc215c822} /* (5, 8, 6) {real, imag} */,
  {32'hc297f78d, 32'h416f8574} /* (5, 8, 5) {real, imag} */,
  {32'h428f4622, 32'hc26ef0dc} /* (5, 8, 4) {real, imag} */,
  {32'h43598d04, 32'h42d0d8be} /* (5, 8, 3) {real, imag} */,
  {32'h431e2e54, 32'hc393dd65} /* (5, 8, 2) {real, imag} */,
  {32'h43281039, 32'h43ccec91} /* (5, 8, 1) {real, imag} */,
  {32'h445a4c22, 32'h00000000} /* (5, 8, 0) {real, imag} */,
  {32'h43a1046c, 32'hc3cfb300} /* (5, 7, 31) {real, imag} */,
  {32'h4332d838, 32'h43c46604} /* (5, 7, 30) {real, imag} */,
  {32'h4371cb39, 32'hc325ae0a} /* (5, 7, 29) {real, imag} */,
  {32'h4209d944, 32'h42d9b7b8} /* (5, 7, 28) {real, imag} */,
  {32'hc2c0b510, 32'h42099a7e} /* (5, 7, 27) {real, imag} */,
  {32'h422b782c, 32'h4326ae66} /* (5, 7, 26) {real, imag} */,
  {32'hc2fa46b7, 32'hc2ee0b30} /* (5, 7, 25) {real, imag} */,
  {32'h42050f72, 32'hc343c275} /* (5, 7, 24) {real, imag} */,
  {32'hc30525f4, 32'h42f47cae} /* (5, 7, 23) {real, imag} */,
  {32'h3f00a1d0, 32'h423dc0d6} /* (5, 7, 22) {real, imag} */,
  {32'h420cab12, 32'hc3334542} /* (5, 7, 21) {real, imag} */,
  {32'hc2b0baad, 32'hc30fff2d} /* (5, 7, 20) {real, imag} */,
  {32'h419a289e, 32'h40ee46b4} /* (5, 7, 19) {real, imag} */,
  {32'h41a2f01c, 32'hc21f7c1e} /* (5, 7, 18) {real, imag} */,
  {32'hc118f62c, 32'h4276c855} /* (5, 7, 17) {real, imag} */,
  {32'h41f4e6e8, 32'h00000000} /* (5, 7, 16) {real, imag} */,
  {32'hc118f62c, 32'hc276c855} /* (5, 7, 15) {real, imag} */,
  {32'h41a2f01c, 32'h421f7c1e} /* (5, 7, 14) {real, imag} */,
  {32'h419a289e, 32'hc0ee46b4} /* (5, 7, 13) {real, imag} */,
  {32'hc2b0baad, 32'h430fff2d} /* (5, 7, 12) {real, imag} */,
  {32'h420cab12, 32'h43334542} /* (5, 7, 11) {real, imag} */,
  {32'h3f00a1d0, 32'hc23dc0d6} /* (5, 7, 10) {real, imag} */,
  {32'hc30525f4, 32'hc2f47cae} /* (5, 7, 9) {real, imag} */,
  {32'h42050f72, 32'h4343c275} /* (5, 7, 8) {real, imag} */,
  {32'hc2fa46b7, 32'h42ee0b30} /* (5, 7, 7) {real, imag} */,
  {32'h422b782c, 32'hc326ae66} /* (5, 7, 6) {real, imag} */,
  {32'hc2c0b510, 32'hc2099a7e} /* (5, 7, 5) {real, imag} */,
  {32'h4209d944, 32'hc2d9b7b8} /* (5, 7, 4) {real, imag} */,
  {32'h4371cb39, 32'h4325ae0a} /* (5, 7, 3) {real, imag} */,
  {32'h4332d838, 32'hc3c46604} /* (5, 7, 2) {real, imag} */,
  {32'h43a1046c, 32'h43cfb300} /* (5, 7, 1) {real, imag} */,
  {32'h448a2d7f, 32'h00000000} /* (5, 7, 0) {real, imag} */,
  {32'h43e8ee86, 32'hc3b65ccc} /* (5, 6, 31) {real, imag} */,
  {32'hc29a4d72, 32'h438d7caa} /* (5, 6, 30) {real, imag} */,
  {32'h434ea4f6, 32'h4201ff35} /* (5, 6, 29) {real, imag} */,
  {32'h428108cf, 32'hc1189688} /* (5, 6, 28) {real, imag} */,
  {32'hc2078244, 32'hc1ce49f8} /* (5, 6, 27) {real, imag} */,
  {32'h42348035, 32'hc1474846} /* (5, 6, 26) {real, imag} */,
  {32'h422e1a76, 32'hc28fc9a2} /* (5, 6, 25) {real, imag} */,
  {32'hc2a613ce, 32'hc13f71e0} /* (5, 6, 24) {real, imag} */,
  {32'hc20afbd6, 32'h4195daa4} /* (5, 6, 23) {real, imag} */,
  {32'hc2689792, 32'hc0d77590} /* (5, 6, 22) {real, imag} */,
  {32'hc29232aa, 32'hc286c9f2} /* (5, 6, 21) {real, imag} */,
  {32'h4231a2f4, 32'h42d8137c} /* (5, 6, 20) {real, imag} */,
  {32'h3fdf67d0, 32'h4262d0f0} /* (5, 6, 19) {real, imag} */,
  {32'h42d567ed, 32'hc046faa8} /* (5, 6, 18) {real, imag} */,
  {32'h4193ac60, 32'h41538f5d} /* (5, 6, 17) {real, imag} */,
  {32'h424795ae, 32'h00000000} /* (5, 6, 16) {real, imag} */,
  {32'h4193ac60, 32'hc1538f5d} /* (5, 6, 15) {real, imag} */,
  {32'h42d567ed, 32'h4046faa8} /* (5, 6, 14) {real, imag} */,
  {32'h3fdf67d0, 32'hc262d0f0} /* (5, 6, 13) {real, imag} */,
  {32'h4231a2f4, 32'hc2d8137c} /* (5, 6, 12) {real, imag} */,
  {32'hc29232aa, 32'h4286c9f2} /* (5, 6, 11) {real, imag} */,
  {32'hc2689792, 32'h40d77590} /* (5, 6, 10) {real, imag} */,
  {32'hc20afbd6, 32'hc195daa4} /* (5, 6, 9) {real, imag} */,
  {32'hc2a613ce, 32'h413f71e0} /* (5, 6, 8) {real, imag} */,
  {32'h422e1a76, 32'h428fc9a2} /* (5, 6, 7) {real, imag} */,
  {32'h42348035, 32'h41474846} /* (5, 6, 6) {real, imag} */,
  {32'hc2078244, 32'h41ce49f8} /* (5, 6, 5) {real, imag} */,
  {32'h428108cf, 32'h41189688} /* (5, 6, 4) {real, imag} */,
  {32'h434ea4f6, 32'hc201ff35} /* (5, 6, 3) {real, imag} */,
  {32'hc29a4d72, 32'hc38d7caa} /* (5, 6, 2) {real, imag} */,
  {32'h43e8ee86, 32'h43b65ccc} /* (5, 6, 1) {real, imag} */,
  {32'h44b265d8, 32'h00000000} /* (5, 6, 0) {real, imag} */,
  {32'h443acd81, 32'hc3b0eedc} /* (5, 5, 31) {real, imag} */,
  {32'hc285272c, 32'h43569a33} /* (5, 5, 30) {real, imag} */,
  {32'h42c2e145, 32'h42d6434f} /* (5, 5, 29) {real, imag} */,
  {32'h41adfdf2, 32'hc2eecb6b} /* (5, 5, 28) {real, imag} */,
  {32'hc144de98, 32'hc2317c31} /* (5, 5, 27) {real, imag} */,
  {32'h4258f4a7, 32'hc27a97ba} /* (5, 5, 26) {real, imag} */,
  {32'h42831162, 32'hc2cd2ba9} /* (5, 5, 25) {real, imag} */,
  {32'hc2a240aa, 32'hc2361174} /* (5, 5, 24) {real, imag} */,
  {32'hc1cb17c6, 32'h4289576d} /* (5, 5, 23) {real, imag} */,
  {32'hc2a04a15, 32'h40acec5c} /* (5, 5, 22) {real, imag} */,
  {32'h41a386cc, 32'h42922ee0} /* (5, 5, 21) {real, imag} */,
  {32'h427a0fba, 32'hc2bcb1a3} /* (5, 5, 20) {real, imag} */,
  {32'h4217d27b, 32'hc236b9ec} /* (5, 5, 19) {real, imag} */,
  {32'h4129a0d7, 32'h42c783a8} /* (5, 5, 18) {real, imag} */,
  {32'hc2e34a46, 32'hc1a6f17a} /* (5, 5, 17) {real, imag} */,
  {32'h41e21306, 32'h00000000} /* (5, 5, 16) {real, imag} */,
  {32'hc2e34a46, 32'h41a6f17a} /* (5, 5, 15) {real, imag} */,
  {32'h4129a0d7, 32'hc2c783a8} /* (5, 5, 14) {real, imag} */,
  {32'h4217d27b, 32'h4236b9ec} /* (5, 5, 13) {real, imag} */,
  {32'h427a0fba, 32'h42bcb1a3} /* (5, 5, 12) {real, imag} */,
  {32'h41a386cc, 32'hc2922ee0} /* (5, 5, 11) {real, imag} */,
  {32'hc2a04a15, 32'hc0acec5c} /* (5, 5, 10) {real, imag} */,
  {32'hc1cb17c6, 32'hc289576d} /* (5, 5, 9) {real, imag} */,
  {32'hc2a240aa, 32'h42361174} /* (5, 5, 8) {real, imag} */,
  {32'h42831162, 32'h42cd2ba9} /* (5, 5, 7) {real, imag} */,
  {32'h4258f4a7, 32'h427a97ba} /* (5, 5, 6) {real, imag} */,
  {32'hc144de98, 32'h42317c31} /* (5, 5, 5) {real, imag} */,
  {32'h41adfdf2, 32'h42eecb6b} /* (5, 5, 4) {real, imag} */,
  {32'h42c2e145, 32'hc2d6434f} /* (5, 5, 3) {real, imag} */,
  {32'hc285272c, 32'hc3569a33} /* (5, 5, 2) {real, imag} */,
  {32'h443acd81, 32'h43b0eedc} /* (5, 5, 1) {real, imag} */,
  {32'h44badec0, 32'h00000000} /* (5, 5, 0) {real, imag} */,
  {32'h444de130, 32'hc3d070e6} /* (5, 4, 31) {real, imag} */,
  {32'hc2aeb34f, 32'h435c89ca} /* (5, 4, 30) {real, imag} */,
  {32'h42fa4546, 32'h420fd9f4} /* (5, 4, 29) {real, imag} */,
  {32'h42876352, 32'hc29157c5} /* (5, 4, 28) {real, imag} */,
  {32'h425d3d18, 32'hc1290778} /* (5, 4, 27) {real, imag} */,
  {32'h42d80742, 32'h4236f9fa} /* (5, 4, 26) {real, imag} */,
  {32'h424be568, 32'hc1aa6278} /* (5, 4, 25) {real, imag} */,
  {32'hc18b9ed6, 32'h42113e32} /* (5, 4, 24) {real, imag} */,
  {32'hc285de98, 32'hc1b5bd50} /* (5, 4, 23) {real, imag} */,
  {32'h42764984, 32'h428f489c} /* (5, 4, 22) {real, imag} */,
  {32'h418f3fea, 32'hc1d878a4} /* (5, 4, 21) {real, imag} */,
  {32'hc263a36c, 32'h4248f64e} /* (5, 4, 20) {real, imag} */,
  {32'h415ed97e, 32'hc158aacc} /* (5, 4, 19) {real, imag} */,
  {32'h42521bc7, 32'hc19dd985} /* (5, 4, 18) {real, imag} */,
  {32'hc14cfb90, 32'hc146690c} /* (5, 4, 17) {real, imag} */,
  {32'h4255d5ba, 32'h00000000} /* (5, 4, 16) {real, imag} */,
  {32'hc14cfb90, 32'h4146690c} /* (5, 4, 15) {real, imag} */,
  {32'h42521bc7, 32'h419dd985} /* (5, 4, 14) {real, imag} */,
  {32'h415ed97e, 32'h4158aacc} /* (5, 4, 13) {real, imag} */,
  {32'hc263a36c, 32'hc248f64e} /* (5, 4, 12) {real, imag} */,
  {32'h418f3fea, 32'h41d878a4} /* (5, 4, 11) {real, imag} */,
  {32'h42764984, 32'hc28f489c} /* (5, 4, 10) {real, imag} */,
  {32'hc285de98, 32'h41b5bd50} /* (5, 4, 9) {real, imag} */,
  {32'hc18b9ed6, 32'hc2113e32} /* (5, 4, 8) {real, imag} */,
  {32'h424be568, 32'h41aa6278} /* (5, 4, 7) {real, imag} */,
  {32'h42d80742, 32'hc236f9fa} /* (5, 4, 6) {real, imag} */,
  {32'h425d3d18, 32'h41290778} /* (5, 4, 5) {real, imag} */,
  {32'h42876352, 32'h429157c5} /* (5, 4, 4) {real, imag} */,
  {32'h42fa4546, 32'hc20fd9f4} /* (5, 4, 3) {real, imag} */,
  {32'hc2aeb34f, 32'hc35c89ca} /* (5, 4, 2) {real, imag} */,
  {32'h444de130, 32'h43d070e6} /* (5, 4, 1) {real, imag} */,
  {32'h44ba11ba, 32'h00000000} /* (5, 4, 0) {real, imag} */,
  {32'h443d98f0, 32'hc40df1a6} /* (5, 3, 31) {real, imag} */,
  {32'hc2760c8e, 32'h42e0c55c} /* (5, 3, 30) {real, imag} */,
  {32'h43016db9, 32'h4198a780} /* (5, 3, 29) {real, imag} */,
  {32'h41cdbb18, 32'h4111d790} /* (5, 3, 28) {real, imag} */,
  {32'h42ef017e, 32'h407e9a60} /* (5, 3, 27) {real, imag} */,
  {32'h42212f0a, 32'hc29ed2e6} /* (5, 3, 26) {real, imag} */,
  {32'h41b168b2, 32'hc1c2fc12} /* (5, 3, 25) {real, imag} */,
  {32'h41a27bb0, 32'h42657d57} /* (5, 3, 24) {real, imag} */,
  {32'h42ca41cc, 32'h42633664} /* (5, 3, 23) {real, imag} */,
  {32'h41e63d28, 32'h42d5faea} /* (5, 3, 22) {real, imag} */,
  {32'hc12837a8, 32'h416e27a6} /* (5, 3, 21) {real, imag} */,
  {32'hc2aaff99, 32'h42b7c2d6} /* (5, 3, 20) {real, imag} */,
  {32'h429d9c62, 32'hc1c1fdaa} /* (5, 3, 19) {real, imag} */,
  {32'h42254693, 32'hc241c987} /* (5, 3, 18) {real, imag} */,
  {32'h4213b1fa, 32'hc1a2796e} /* (5, 3, 17) {real, imag} */,
  {32'hc1ebcfa5, 32'h00000000} /* (5, 3, 16) {real, imag} */,
  {32'h4213b1fa, 32'h41a2796e} /* (5, 3, 15) {real, imag} */,
  {32'h42254693, 32'h4241c987} /* (5, 3, 14) {real, imag} */,
  {32'h429d9c62, 32'h41c1fdaa} /* (5, 3, 13) {real, imag} */,
  {32'hc2aaff99, 32'hc2b7c2d6} /* (5, 3, 12) {real, imag} */,
  {32'hc12837a8, 32'hc16e27a6} /* (5, 3, 11) {real, imag} */,
  {32'h41e63d28, 32'hc2d5faea} /* (5, 3, 10) {real, imag} */,
  {32'h42ca41cc, 32'hc2633664} /* (5, 3, 9) {real, imag} */,
  {32'h41a27bb0, 32'hc2657d57} /* (5, 3, 8) {real, imag} */,
  {32'h41b168b2, 32'h41c2fc12} /* (5, 3, 7) {real, imag} */,
  {32'h42212f0a, 32'h429ed2e6} /* (5, 3, 6) {real, imag} */,
  {32'h42ef017e, 32'hc07e9a60} /* (5, 3, 5) {real, imag} */,
  {32'h41cdbb18, 32'hc111d790} /* (5, 3, 4) {real, imag} */,
  {32'h43016db9, 32'hc198a780} /* (5, 3, 3) {real, imag} */,
  {32'hc2760c8e, 32'hc2e0c55c} /* (5, 3, 2) {real, imag} */,
  {32'h443d98f0, 32'h440df1a6} /* (5, 3, 1) {real, imag} */,
  {32'h44cae2c5, 32'h00000000} /* (5, 3, 0) {real, imag} */,
  {32'h443510cd, 32'hc403ee29} /* (5, 2, 31) {real, imag} */,
  {32'hc1144cc8, 32'hc1d9fa8e} /* (5, 2, 30) {real, imag} */,
  {32'h42d9adba, 32'h424ae05d} /* (5, 2, 29) {real, imag} */,
  {32'h42125e2e, 32'hc2b58bb0} /* (5, 2, 28) {real, imag} */,
  {32'h4277e9f9, 32'h401a2360} /* (5, 2, 27) {real, imag} */,
  {32'hc0a57e14, 32'hc22621fa} /* (5, 2, 26) {real, imag} */,
  {32'hc3149383, 32'hc2a2afdf} /* (5, 2, 25) {real, imag} */,
  {32'hc2340a56, 32'hc2069033} /* (5, 2, 24) {real, imag} */,
  {32'hc28e1727, 32'h4241c4e8} /* (5, 2, 23) {real, imag} */,
  {32'hc283b5d3, 32'hc2994ff9} /* (5, 2, 22) {real, imag} */,
  {32'h40be91f0, 32'h4296cb9d} /* (5, 2, 21) {real, imag} */,
  {32'h41adb6c9, 32'hc0c77b54} /* (5, 2, 20) {real, imag} */,
  {32'hc1adb9ec, 32'hc2095f72} /* (5, 2, 19) {real, imag} */,
  {32'hc1c3b983, 32'hc241b902} /* (5, 2, 18) {real, imag} */,
  {32'h4123fac3, 32'h4299dc32} /* (5, 2, 17) {real, imag} */,
  {32'hc1c7ac14, 32'h00000000} /* (5, 2, 16) {real, imag} */,
  {32'h4123fac3, 32'hc299dc32} /* (5, 2, 15) {real, imag} */,
  {32'hc1c3b983, 32'h4241b902} /* (5, 2, 14) {real, imag} */,
  {32'hc1adb9ec, 32'h42095f72} /* (5, 2, 13) {real, imag} */,
  {32'h41adb6c9, 32'h40c77b54} /* (5, 2, 12) {real, imag} */,
  {32'h40be91f0, 32'hc296cb9d} /* (5, 2, 11) {real, imag} */,
  {32'hc283b5d3, 32'h42994ff9} /* (5, 2, 10) {real, imag} */,
  {32'hc28e1727, 32'hc241c4e8} /* (5, 2, 9) {real, imag} */,
  {32'hc2340a56, 32'h42069033} /* (5, 2, 8) {real, imag} */,
  {32'hc3149383, 32'h42a2afdf} /* (5, 2, 7) {real, imag} */,
  {32'hc0a57e14, 32'h422621fa} /* (5, 2, 6) {real, imag} */,
  {32'h4277e9f9, 32'hc01a2360} /* (5, 2, 5) {real, imag} */,
  {32'h42125e2e, 32'h42b58bb0} /* (5, 2, 4) {real, imag} */,
  {32'h42d9adba, 32'hc24ae05d} /* (5, 2, 3) {real, imag} */,
  {32'hc1144cc8, 32'h41d9fa8e} /* (5, 2, 2) {real, imag} */,
  {32'h443510cd, 32'h4403ee29} /* (5, 2, 1) {real, imag} */,
  {32'h44e66f2d, 32'h00000000} /* (5, 2, 0) {real, imag} */,
  {32'h4447ae08, 32'hc3cff9b3} /* (5, 1, 31) {real, imag} */,
  {32'hc22687e8, 32'hc32823a8} /* (5, 1, 30) {real, imag} */,
  {32'h42e3e257, 32'hc13059b8} /* (5, 1, 29) {real, imag} */,
  {32'h42b95bb3, 32'hc30098bb} /* (5, 1, 28) {real, imag} */,
  {32'hc2c577b0, 32'h4212f376} /* (5, 1, 27) {real, imag} */,
  {32'hc24932c2, 32'hc180c422} /* (5, 1, 26) {real, imag} */,
  {32'hc24dee94, 32'h43324262} /* (5, 1, 25) {real, imag} */,
  {32'h42e23ebe, 32'hc2ddcae6} /* (5, 1, 24) {real, imag} */,
  {32'hc1c486f9, 32'hc1f03f2a} /* (5, 1, 23) {real, imag} */,
  {32'hc10db809, 32'h4214cb33} /* (5, 1, 22) {real, imag} */,
  {32'hc1a2ff4a, 32'h411d2e88} /* (5, 1, 21) {real, imag} */,
  {32'h4240ed93, 32'h41ba28e3} /* (5, 1, 20) {real, imag} */,
  {32'hc2bf42ec, 32'hc22760bc} /* (5, 1, 19) {real, imag} */,
  {32'h41d94afa, 32'hc1322920} /* (5, 1, 18) {real, imag} */,
  {32'h3ecf1e80, 32'hc2298f90} /* (5, 1, 17) {real, imag} */,
  {32'hbf1db480, 32'h00000000} /* (5, 1, 16) {real, imag} */,
  {32'h3ecf1e80, 32'h42298f90} /* (5, 1, 15) {real, imag} */,
  {32'h41d94afa, 32'h41322920} /* (5, 1, 14) {real, imag} */,
  {32'hc2bf42ec, 32'h422760bc} /* (5, 1, 13) {real, imag} */,
  {32'h4240ed93, 32'hc1ba28e3} /* (5, 1, 12) {real, imag} */,
  {32'hc1a2ff4a, 32'hc11d2e88} /* (5, 1, 11) {real, imag} */,
  {32'hc10db809, 32'hc214cb33} /* (5, 1, 10) {real, imag} */,
  {32'hc1c486f9, 32'h41f03f2a} /* (5, 1, 9) {real, imag} */,
  {32'h42e23ebe, 32'h42ddcae6} /* (5, 1, 8) {real, imag} */,
  {32'hc24dee94, 32'hc3324262} /* (5, 1, 7) {real, imag} */,
  {32'hc24932c2, 32'h4180c422} /* (5, 1, 6) {real, imag} */,
  {32'hc2c577b0, 32'hc212f376} /* (5, 1, 5) {real, imag} */,
  {32'h42b95bb3, 32'h430098bb} /* (5, 1, 4) {real, imag} */,
  {32'h42e3e257, 32'h413059b8} /* (5, 1, 3) {real, imag} */,
  {32'hc22687e8, 32'h432823a8} /* (5, 1, 2) {real, imag} */,
  {32'h4447ae08, 32'h43cff9b3} /* (5, 1, 1) {real, imag} */,
  {32'h44f4a426, 32'h00000000} /* (5, 1, 0) {real, imag} */,
  {32'h44588a52, 32'hc415dae1} /* (5, 0, 31) {real, imag} */,
  {32'h4247967e, 32'hc2dee23e} /* (5, 0, 30) {real, imag} */,
  {32'h42dbe5ac, 32'h4254ffaa} /* (5, 0, 29) {real, imag} */,
  {32'hc1829b56, 32'hc271b0d3} /* (5, 0, 28) {real, imag} */,
  {32'hc25c5a1a, 32'hc14b4642} /* (5, 0, 27) {real, imag} */,
  {32'hc2808254, 32'h41c186e0} /* (5, 0, 26) {real, imag} */,
  {32'hc23a297c, 32'h42176e5c} /* (5, 0, 25) {real, imag} */,
  {32'h424f1056, 32'hc0dab984} /* (5, 0, 24) {real, imag} */,
  {32'hc1b7f0aa, 32'hc22024ca} /* (5, 0, 23) {real, imag} */,
  {32'hc1f10ab8, 32'h4116f3a0} /* (5, 0, 22) {real, imag} */,
  {32'hc0ef6838, 32'hc1e02a70} /* (5, 0, 21) {real, imag} */,
  {32'h41f3265e, 32'h4205f818} /* (5, 0, 20) {real, imag} */,
  {32'h41e67428, 32'hc17cbddc} /* (5, 0, 19) {real, imag} */,
  {32'hc1b83a43, 32'h429c8bae} /* (5, 0, 18) {real, imag} */,
  {32'hc210932f, 32'hc17796f4} /* (5, 0, 17) {real, imag} */,
  {32'h4224425a, 32'h00000000} /* (5, 0, 16) {real, imag} */,
  {32'hc210932f, 32'h417796f4} /* (5, 0, 15) {real, imag} */,
  {32'hc1b83a43, 32'hc29c8bae} /* (5, 0, 14) {real, imag} */,
  {32'h41e67428, 32'h417cbddc} /* (5, 0, 13) {real, imag} */,
  {32'h41f3265e, 32'hc205f818} /* (5, 0, 12) {real, imag} */,
  {32'hc0ef6838, 32'h41e02a70} /* (5, 0, 11) {real, imag} */,
  {32'hc1f10ab8, 32'hc116f3a0} /* (5, 0, 10) {real, imag} */,
  {32'hc1b7f0aa, 32'h422024ca} /* (5, 0, 9) {real, imag} */,
  {32'h424f1056, 32'h40dab984} /* (5, 0, 8) {real, imag} */,
  {32'hc23a297c, 32'hc2176e5c} /* (5, 0, 7) {real, imag} */,
  {32'hc2808254, 32'hc1c186e0} /* (5, 0, 6) {real, imag} */,
  {32'hc25c5a1a, 32'h414b4642} /* (5, 0, 5) {real, imag} */,
  {32'hc1829b56, 32'h4271b0d3} /* (5, 0, 4) {real, imag} */,
  {32'h42dbe5ac, 32'hc254ffaa} /* (5, 0, 3) {real, imag} */,
  {32'h4247967e, 32'h42dee23e} /* (5, 0, 2) {real, imag} */,
  {32'h44588a52, 32'h4415dae1} /* (5, 0, 1) {real, imag} */,
  {32'h450283e6, 32'h00000000} /* (5, 0, 0) {real, imag} */,
  {32'hc3462a88, 32'h426d6720} /* (4, 31, 31) {real, imag} */,
  {32'h43d0de82, 32'hc2f61456} /* (4, 31, 30) {real, imag} */,
  {32'h4336da98, 32'hc259bc15} /* (4, 31, 29) {real, imag} */,
  {32'hc2f4ef42, 32'hc2ab94b8} /* (4, 31, 28) {real, imag} */,
  {32'h4257e92e, 32'hc15c5690} /* (4, 31, 27) {real, imag} */,
  {32'hc28e6c5e, 32'h429d11ed} /* (4, 31, 26) {real, imag} */,
  {32'hc0da0330, 32'hc1f10099} /* (4, 31, 25) {real, imag} */,
  {32'h4252be99, 32'h4189823a} /* (4, 31, 24) {real, imag} */,
  {32'hc20eb817, 32'h4249b103} /* (4, 31, 23) {real, imag} */,
  {32'h42142641, 32'h42076d31} /* (4, 31, 22) {real, imag} */,
  {32'hc20e0c79, 32'hc22d8768} /* (4, 31, 21) {real, imag} */,
  {32'hc2026823, 32'h40372724} /* (4, 31, 20) {real, imag} */,
  {32'h41bcfbba, 32'h4201d45a} /* (4, 31, 19) {real, imag} */,
  {32'h40f70dac, 32'hc205e93a} /* (4, 31, 18) {real, imag} */,
  {32'h4222f756, 32'hc1afa3a4} /* (4, 31, 17) {real, imag} */,
  {32'hc2b0f278, 32'h00000000} /* (4, 31, 16) {real, imag} */,
  {32'h4222f756, 32'h41afa3a4} /* (4, 31, 15) {real, imag} */,
  {32'h40f70dac, 32'h4205e93a} /* (4, 31, 14) {real, imag} */,
  {32'h41bcfbba, 32'hc201d45a} /* (4, 31, 13) {real, imag} */,
  {32'hc2026823, 32'hc0372724} /* (4, 31, 12) {real, imag} */,
  {32'hc20e0c79, 32'h422d8768} /* (4, 31, 11) {real, imag} */,
  {32'h42142641, 32'hc2076d31} /* (4, 31, 10) {real, imag} */,
  {32'hc20eb817, 32'hc249b103} /* (4, 31, 9) {real, imag} */,
  {32'h4252be99, 32'hc189823a} /* (4, 31, 8) {real, imag} */,
  {32'hc0da0330, 32'h41f10099} /* (4, 31, 7) {real, imag} */,
  {32'hc28e6c5e, 32'hc29d11ed} /* (4, 31, 6) {real, imag} */,
  {32'h4257e92e, 32'h415c5690} /* (4, 31, 5) {real, imag} */,
  {32'hc2f4ef42, 32'h42ab94b8} /* (4, 31, 4) {real, imag} */,
  {32'h4336da98, 32'h4259bc15} /* (4, 31, 3) {real, imag} */,
  {32'h43d0de82, 32'h42f61456} /* (4, 31, 2) {real, imag} */,
  {32'hc3462a88, 32'hc26d6720} /* (4, 31, 1) {real, imag} */,
  {32'h44604fbc, 32'h00000000} /* (4, 31, 0) {real, imag} */,
  {32'hc408da75, 32'h420f6070} /* (4, 30, 31) {real, imag} */,
  {32'h4420cc7e, 32'hc309d191} /* (4, 30, 30) {real, imag} */,
  {32'h433e44fe, 32'hc200241b} /* (4, 30, 29) {real, imag} */,
  {32'hc31e7236, 32'h41099b60} /* (4, 30, 28) {real, imag} */,
  {32'h4264081c, 32'hc1f3c99c} /* (4, 30, 27) {real, imag} */,
  {32'hc26bc67e, 32'h429b5ad9} /* (4, 30, 26) {real, imag} */,
  {32'hc14b14dc, 32'h40827d78} /* (4, 30, 25) {real, imag} */,
  {32'h42a8abf4, 32'hc1c0572a} /* (4, 30, 24) {real, imag} */,
  {32'h41acdc7a, 32'h4187b744} /* (4, 30, 23) {real, imag} */,
  {32'h40666990, 32'hc245cfd5} /* (4, 30, 22) {real, imag} */,
  {32'h40fa0d9c, 32'hc2283ea4} /* (4, 30, 21) {real, imag} */,
  {32'h420b5665, 32'hc0c355c2} /* (4, 30, 20) {real, imag} */,
  {32'h41d78d36, 32'hc101ea58} /* (4, 30, 19) {real, imag} */,
  {32'hc1ed353e, 32'hc29ef0de} /* (4, 30, 18) {real, imag} */,
  {32'h423ee5f5, 32'hc20ba779} /* (4, 30, 17) {real, imag} */,
  {32'hc26e71d4, 32'h00000000} /* (4, 30, 16) {real, imag} */,
  {32'h423ee5f5, 32'h420ba779} /* (4, 30, 15) {real, imag} */,
  {32'hc1ed353e, 32'h429ef0de} /* (4, 30, 14) {real, imag} */,
  {32'h41d78d36, 32'h4101ea58} /* (4, 30, 13) {real, imag} */,
  {32'h420b5665, 32'h40c355c2} /* (4, 30, 12) {real, imag} */,
  {32'h40fa0d9c, 32'h42283ea4} /* (4, 30, 11) {real, imag} */,
  {32'h40666990, 32'h4245cfd5} /* (4, 30, 10) {real, imag} */,
  {32'h41acdc7a, 32'hc187b744} /* (4, 30, 9) {real, imag} */,
  {32'h42a8abf4, 32'h41c0572a} /* (4, 30, 8) {real, imag} */,
  {32'hc14b14dc, 32'hc0827d78} /* (4, 30, 7) {real, imag} */,
  {32'hc26bc67e, 32'hc29b5ad9} /* (4, 30, 6) {real, imag} */,
  {32'h4264081c, 32'h41f3c99c} /* (4, 30, 5) {real, imag} */,
  {32'hc31e7236, 32'hc1099b60} /* (4, 30, 4) {real, imag} */,
  {32'h433e44fe, 32'h4200241b} /* (4, 30, 3) {real, imag} */,
  {32'h4420cc7e, 32'h4309d191} /* (4, 30, 2) {real, imag} */,
  {32'hc408da75, 32'hc20f6070} /* (4, 30, 1) {real, imag} */,
  {32'h442b6bb4, 32'h00000000} /* (4, 30, 0) {real, imag} */,
  {32'hc42d4510, 32'hc10d4000} /* (4, 29, 31) {real, imag} */,
  {32'h443ec81d, 32'hc256a988} /* (4, 29, 30) {real, imag} */,
  {32'hc0021490, 32'hc1fe2773} /* (4, 29, 29) {real, imag} */,
  {32'hc30f596a, 32'h42c1da0c} /* (4, 29, 28) {real, imag} */,
  {32'h4281ba64, 32'h40821e50} /* (4, 29, 27) {real, imag} */,
  {32'h428e12f7, 32'h42b5d56d} /* (4, 29, 26) {real, imag} */,
  {32'hc30abc5b, 32'hc10e8728} /* (4, 29, 25) {real, imag} */,
  {32'h42f33dab, 32'hc2cb9e28} /* (4, 29, 24) {real, imag} */,
  {32'hc28d6100, 32'hc21c4afc} /* (4, 29, 23) {real, imag} */,
  {32'hc21512df, 32'hc2cdff92} /* (4, 29, 22) {real, imag} */,
  {32'h41f592e9, 32'hc2c15568} /* (4, 29, 21) {real, imag} */,
  {32'h42299c19, 32'h42beb600} /* (4, 29, 20) {real, imag} */,
  {32'hc192d030, 32'hc2576a9b} /* (4, 29, 19) {real, imag} */,
  {32'hc225e483, 32'hc1e62835} /* (4, 29, 18) {real, imag} */,
  {32'h41ccf21a, 32'hc0a1d1b0} /* (4, 29, 17) {real, imag} */,
  {32'hc249a9ae, 32'h00000000} /* (4, 29, 16) {real, imag} */,
  {32'h41ccf21a, 32'h40a1d1b0} /* (4, 29, 15) {real, imag} */,
  {32'hc225e483, 32'h41e62835} /* (4, 29, 14) {real, imag} */,
  {32'hc192d030, 32'h42576a9b} /* (4, 29, 13) {real, imag} */,
  {32'h42299c19, 32'hc2beb600} /* (4, 29, 12) {real, imag} */,
  {32'h41f592e9, 32'h42c15568} /* (4, 29, 11) {real, imag} */,
  {32'hc21512df, 32'h42cdff92} /* (4, 29, 10) {real, imag} */,
  {32'hc28d6100, 32'h421c4afc} /* (4, 29, 9) {real, imag} */,
  {32'h42f33dab, 32'h42cb9e28} /* (4, 29, 8) {real, imag} */,
  {32'hc30abc5b, 32'h410e8728} /* (4, 29, 7) {real, imag} */,
  {32'h428e12f7, 32'hc2b5d56d} /* (4, 29, 6) {real, imag} */,
  {32'h4281ba64, 32'hc0821e50} /* (4, 29, 5) {real, imag} */,
  {32'hc30f596a, 32'hc2c1da0c} /* (4, 29, 4) {real, imag} */,
  {32'hc0021490, 32'h41fe2773} /* (4, 29, 3) {real, imag} */,
  {32'h443ec81d, 32'h4256a988} /* (4, 29, 2) {real, imag} */,
  {32'hc42d4510, 32'h410d4000} /* (4, 29, 1) {real, imag} */,
  {32'h4414e045, 32'h00000000} /* (4, 29, 0) {real, imag} */,
  {32'hc4392fd3, 32'hc14bcda0} /* (4, 28, 31) {real, imag} */,
  {32'h44195331, 32'hc0b7d420} /* (4, 28, 30) {real, imag} */,
  {32'h435c82e5, 32'hc2b4552e} /* (4, 28, 29) {real, imag} */,
  {32'hc364ab64, 32'h41977520} /* (4, 28, 28) {real, imag} */,
  {32'h433492a4, 32'hc28f18fe} /* (4, 28, 27) {real, imag} */,
  {32'h4345f3d7, 32'h416e8312} /* (4, 28, 26) {real, imag} */,
  {32'hc2d9fdb0, 32'h4209a34a} /* (4, 28, 25) {real, imag} */,
  {32'h423ada98, 32'hc2aa3d09} /* (4, 28, 24) {real, imag} */,
  {32'h417c0fd4, 32'hc2be40ee} /* (4, 28, 23) {real, imag} */,
  {32'hc1e44111, 32'h42086372} /* (4, 28, 22) {real, imag} */,
  {32'hc2da4696, 32'hc2534596} /* (4, 28, 21) {real, imag} */,
  {32'hbfb8f768, 32'hc174b74a} /* (4, 28, 20) {real, imag} */,
  {32'hc1d5939d, 32'h422f1f40} /* (4, 28, 19) {real, imag} */,
  {32'h41d7f64c, 32'h41c0a91b} /* (4, 28, 18) {real, imag} */,
  {32'h42179692, 32'h41d50e6f} /* (4, 28, 17) {real, imag} */,
  {32'hc237cac8, 32'h00000000} /* (4, 28, 16) {real, imag} */,
  {32'h42179692, 32'hc1d50e6f} /* (4, 28, 15) {real, imag} */,
  {32'h41d7f64c, 32'hc1c0a91b} /* (4, 28, 14) {real, imag} */,
  {32'hc1d5939d, 32'hc22f1f40} /* (4, 28, 13) {real, imag} */,
  {32'hbfb8f768, 32'h4174b74a} /* (4, 28, 12) {real, imag} */,
  {32'hc2da4696, 32'h42534596} /* (4, 28, 11) {real, imag} */,
  {32'hc1e44111, 32'hc2086372} /* (4, 28, 10) {real, imag} */,
  {32'h417c0fd4, 32'h42be40ee} /* (4, 28, 9) {real, imag} */,
  {32'h423ada98, 32'h42aa3d09} /* (4, 28, 8) {real, imag} */,
  {32'hc2d9fdb0, 32'hc209a34a} /* (4, 28, 7) {real, imag} */,
  {32'h4345f3d7, 32'hc16e8312} /* (4, 28, 6) {real, imag} */,
  {32'h433492a4, 32'h428f18fe} /* (4, 28, 5) {real, imag} */,
  {32'hc364ab64, 32'hc1977520} /* (4, 28, 4) {real, imag} */,
  {32'h435c82e5, 32'h42b4552e} /* (4, 28, 3) {real, imag} */,
  {32'h44195331, 32'h40b7d420} /* (4, 28, 2) {real, imag} */,
  {32'hc4392fd3, 32'h414bcda0} /* (4, 28, 1) {real, imag} */,
  {32'h4415f723, 32'h00000000} /* (4, 28, 0) {real, imag} */,
  {32'hc465b10a, 32'h42f4f6bc} /* (4, 27, 31) {real, imag} */,
  {32'h442ce203, 32'hc0dc9e98} /* (4, 27, 30) {real, imag} */,
  {32'h42d116a1, 32'hc300afc9} /* (4, 27, 29) {real, imag} */,
  {32'hc38944b9, 32'h41e6429c} /* (4, 27, 28) {real, imag} */,
  {32'h431eb158, 32'hc2daf0db} /* (4, 27, 27) {real, imag} */,
  {32'h411d0288, 32'hc22cce7c} /* (4, 27, 26) {real, imag} */,
  {32'hc284a832, 32'h41ecd8e5} /* (4, 27, 25) {real, imag} */,
  {32'h424f8078, 32'hc318b16e} /* (4, 27, 24) {real, imag} */,
  {32'h41936bba, 32'h4305d34e} /* (4, 27, 23) {real, imag} */,
  {32'hc27df722, 32'h421a51c8} /* (4, 27, 22) {real, imag} */,
  {32'h42d43f5a, 32'hc22b54b6} /* (4, 27, 21) {real, imag} */,
  {32'hc2f4ae96, 32'hc2f2202e} /* (4, 27, 20) {real, imag} */,
  {32'h418151ca, 32'h418d0061} /* (4, 27, 19) {real, imag} */,
  {32'h419abde8, 32'hc301a751} /* (4, 27, 18) {real, imag} */,
  {32'hc0e01b09, 32'h41c16c3f} /* (4, 27, 17) {real, imag} */,
  {32'hc2b94ad5, 32'h00000000} /* (4, 27, 16) {real, imag} */,
  {32'hc0e01b09, 32'hc1c16c3f} /* (4, 27, 15) {real, imag} */,
  {32'h419abde8, 32'h4301a751} /* (4, 27, 14) {real, imag} */,
  {32'h418151ca, 32'hc18d0061} /* (4, 27, 13) {real, imag} */,
  {32'hc2f4ae96, 32'h42f2202e} /* (4, 27, 12) {real, imag} */,
  {32'h42d43f5a, 32'h422b54b6} /* (4, 27, 11) {real, imag} */,
  {32'hc27df722, 32'hc21a51c8} /* (4, 27, 10) {real, imag} */,
  {32'h41936bba, 32'hc305d34e} /* (4, 27, 9) {real, imag} */,
  {32'h424f8078, 32'h4318b16e} /* (4, 27, 8) {real, imag} */,
  {32'hc284a832, 32'hc1ecd8e5} /* (4, 27, 7) {real, imag} */,
  {32'h411d0288, 32'h422cce7c} /* (4, 27, 6) {real, imag} */,
  {32'h431eb158, 32'h42daf0db} /* (4, 27, 5) {real, imag} */,
  {32'hc38944b9, 32'hc1e6429c} /* (4, 27, 4) {real, imag} */,
  {32'h42d116a1, 32'h4300afc9} /* (4, 27, 3) {real, imag} */,
  {32'h442ce203, 32'h40dc9e98} /* (4, 27, 2) {real, imag} */,
  {32'hc465b10a, 32'hc2f4f6bc} /* (4, 27, 1) {real, imag} */,
  {32'h441c03cc, 32'h00000000} /* (4, 27, 0) {real, imag} */,
  {32'hc462ec6f, 32'h436ec5dc} /* (4, 26, 31) {real, imag} */,
  {32'h443bf48b, 32'hc22d2816} /* (4, 26, 30) {real, imag} */,
  {32'hc14a50d0, 32'hc2f9923c} /* (4, 26, 29) {real, imag} */,
  {32'hc33783dc, 32'hc1f1be06} /* (4, 26, 28) {real, imag} */,
  {32'h4329ee63, 32'h42065bd1} /* (4, 26, 27) {real, imag} */,
  {32'h42685516, 32'h40e2870c} /* (4, 26, 26) {real, imag} */,
  {32'hc15fcfbc, 32'hc205b5d0} /* (4, 26, 25) {real, imag} */,
  {32'h40e9d858, 32'hc28cac05} /* (4, 26, 24) {real, imag} */,
  {32'h4299c794, 32'hbfbb3500} /* (4, 26, 23) {real, imag} */,
  {32'hc1c5fe6e, 32'hc24284bb} /* (4, 26, 22) {real, imag} */,
  {32'h42301782, 32'hc1e49f20} /* (4, 26, 21) {real, imag} */,
  {32'hc1c83206, 32'h426ead7c} /* (4, 26, 20) {real, imag} */,
  {32'h42a31692, 32'hc17beacc} /* (4, 26, 19) {real, imag} */,
  {32'hc13a6a10, 32'h41b2126e} /* (4, 26, 18) {real, imag} */,
  {32'hc20e634c, 32'hc212ab48} /* (4, 26, 17) {real, imag} */,
  {32'hc203d2b2, 32'h00000000} /* (4, 26, 16) {real, imag} */,
  {32'hc20e634c, 32'h4212ab48} /* (4, 26, 15) {real, imag} */,
  {32'hc13a6a10, 32'hc1b2126e} /* (4, 26, 14) {real, imag} */,
  {32'h42a31692, 32'h417beacc} /* (4, 26, 13) {real, imag} */,
  {32'hc1c83206, 32'hc26ead7c} /* (4, 26, 12) {real, imag} */,
  {32'h42301782, 32'h41e49f20} /* (4, 26, 11) {real, imag} */,
  {32'hc1c5fe6e, 32'h424284bb} /* (4, 26, 10) {real, imag} */,
  {32'h4299c794, 32'h3fbb3500} /* (4, 26, 9) {real, imag} */,
  {32'h40e9d858, 32'h428cac05} /* (4, 26, 8) {real, imag} */,
  {32'hc15fcfbc, 32'h4205b5d0} /* (4, 26, 7) {real, imag} */,
  {32'h42685516, 32'hc0e2870c} /* (4, 26, 6) {real, imag} */,
  {32'h4329ee63, 32'hc2065bd1} /* (4, 26, 5) {real, imag} */,
  {32'hc33783dc, 32'h41f1be06} /* (4, 26, 4) {real, imag} */,
  {32'hc14a50d0, 32'h42f9923c} /* (4, 26, 3) {real, imag} */,
  {32'h443bf48b, 32'h422d2816} /* (4, 26, 2) {real, imag} */,
  {32'hc462ec6f, 32'hc36ec5dc} /* (4, 26, 1) {real, imag} */,
  {32'h4404ff53, 32'h00000000} /* (4, 26, 0) {real, imag} */,
  {32'hc4886cd2, 32'h43291975} /* (4, 25, 31) {real, imag} */,
  {32'h443f5c10, 32'hc1cc2802} /* (4, 25, 30) {real, imag} */,
  {32'h42c74ce9, 32'hc329170c} /* (4, 25, 29) {real, imag} */,
  {32'hc33182b2, 32'h42878efb} /* (4, 25, 28) {real, imag} */,
  {32'h43329900, 32'hc21677ad} /* (4, 25, 27) {real, imag} */,
  {32'h419b335a, 32'hc19cbfda} /* (4, 25, 26) {real, imag} */,
  {32'hc25cba1d, 32'h42f696da} /* (4, 25, 25) {real, imag} */,
  {32'h4254f288, 32'hc2eb1740} /* (4, 25, 24) {real, imag} */,
  {32'hc1327bbe, 32'hc2b9ef54} /* (4, 25, 23) {real, imag} */,
  {32'h42ca71ef, 32'h4297929c} /* (4, 25, 22) {real, imag} */,
  {32'h42a98b9e, 32'h4206abfe} /* (4, 25, 21) {real, imag} */,
  {32'hc0f68fc8, 32'h4249bc93} /* (4, 25, 20) {real, imag} */,
  {32'hc26105da, 32'h4182c408} /* (4, 25, 19) {real, imag} */,
  {32'hc2425f03, 32'hc2c3e443} /* (4, 25, 18) {real, imag} */,
  {32'h41fbd412, 32'h42e9507e} /* (4, 25, 17) {real, imag} */,
  {32'hc2428e09, 32'h00000000} /* (4, 25, 16) {real, imag} */,
  {32'h41fbd412, 32'hc2e9507e} /* (4, 25, 15) {real, imag} */,
  {32'hc2425f03, 32'h42c3e443} /* (4, 25, 14) {real, imag} */,
  {32'hc26105da, 32'hc182c408} /* (4, 25, 13) {real, imag} */,
  {32'hc0f68fc8, 32'hc249bc93} /* (4, 25, 12) {real, imag} */,
  {32'h42a98b9e, 32'hc206abfe} /* (4, 25, 11) {real, imag} */,
  {32'h42ca71ef, 32'hc297929c} /* (4, 25, 10) {real, imag} */,
  {32'hc1327bbe, 32'h42b9ef54} /* (4, 25, 9) {real, imag} */,
  {32'h4254f288, 32'h42eb1740} /* (4, 25, 8) {real, imag} */,
  {32'hc25cba1d, 32'hc2f696da} /* (4, 25, 7) {real, imag} */,
  {32'h419b335a, 32'h419cbfda} /* (4, 25, 6) {real, imag} */,
  {32'h43329900, 32'h421677ad} /* (4, 25, 5) {real, imag} */,
  {32'hc33182b2, 32'hc2878efb} /* (4, 25, 4) {real, imag} */,
  {32'h42c74ce9, 32'h4329170c} /* (4, 25, 3) {real, imag} */,
  {32'h443f5c10, 32'h41cc2802} /* (4, 25, 2) {real, imag} */,
  {32'hc4886cd2, 32'hc3291975} /* (4, 25, 1) {real, imag} */,
  {32'h42c7aa7c, 32'h00000000} /* (4, 25, 0) {real, imag} */,
  {32'hc4a3aaa8, 32'h42b010a2} /* (4, 24, 31) {real, imag} */,
  {32'h44294120, 32'h4304c7b0} /* (4, 24, 30) {real, imag} */,
  {32'hc2239084, 32'hc2b9b1aa} /* (4, 24, 29) {real, imag} */,
  {32'hc3324164, 32'hc198199f} /* (4, 24, 28) {real, imag} */,
  {32'h43144038, 32'hc2eda0a9} /* (4, 24, 27) {real, imag} */,
  {32'hc1add771, 32'hc2efaa1c} /* (4, 24, 26) {real, imag} */,
  {32'hc0d1be08, 32'h410f6804} /* (4, 24, 25) {real, imag} */,
  {32'h42b4890d, 32'hc35da5fa} /* (4, 24, 24) {real, imag} */,
  {32'h416b19fc, 32'hc2130f11} /* (4, 24, 23) {real, imag} */,
  {32'hc0acc850, 32'hc1f96dbb} /* (4, 24, 22) {real, imag} */,
  {32'h4166322a, 32'h4050cce0} /* (4, 24, 21) {real, imag} */,
  {32'hc1687d58, 32'h41cb7940} /* (4, 24, 20) {real, imag} */,
  {32'h41e51a39, 32'h42108554} /* (4, 24, 19) {real, imag} */,
  {32'h41f2d7e8, 32'hc29e4d73} /* (4, 24, 18) {real, imag} */,
  {32'hc1e0c3b4, 32'h429c2f1a} /* (4, 24, 17) {real, imag} */,
  {32'hc2595b63, 32'h00000000} /* (4, 24, 16) {real, imag} */,
  {32'hc1e0c3b4, 32'hc29c2f1a} /* (4, 24, 15) {real, imag} */,
  {32'h41f2d7e8, 32'h429e4d73} /* (4, 24, 14) {real, imag} */,
  {32'h41e51a39, 32'hc2108554} /* (4, 24, 13) {real, imag} */,
  {32'hc1687d58, 32'hc1cb7940} /* (4, 24, 12) {real, imag} */,
  {32'h4166322a, 32'hc050cce0} /* (4, 24, 11) {real, imag} */,
  {32'hc0acc850, 32'h41f96dbb} /* (4, 24, 10) {real, imag} */,
  {32'h416b19fc, 32'h42130f11} /* (4, 24, 9) {real, imag} */,
  {32'h42b4890d, 32'h435da5fa} /* (4, 24, 8) {real, imag} */,
  {32'hc0d1be08, 32'hc10f6804} /* (4, 24, 7) {real, imag} */,
  {32'hc1add771, 32'h42efaa1c} /* (4, 24, 6) {real, imag} */,
  {32'h43144038, 32'h42eda0a9} /* (4, 24, 5) {real, imag} */,
  {32'hc3324164, 32'h4198199f} /* (4, 24, 4) {real, imag} */,
  {32'hc2239084, 32'h42b9b1aa} /* (4, 24, 3) {real, imag} */,
  {32'h44294120, 32'hc304c7b0} /* (4, 24, 2) {real, imag} */,
  {32'hc4a3aaa8, 32'hc2b010a2} /* (4, 24, 1) {real, imag} */,
  {32'h436934f6, 32'h00000000} /* (4, 24, 0) {real, imag} */,
  {32'hc4a0d6b7, 32'hc20453f8} /* (4, 23, 31) {real, imag} */,
  {32'h44236956, 32'h43493776} /* (4, 23, 30) {real, imag} */,
  {32'hc240485c, 32'hc1d9cc42} /* (4, 23, 29) {real, imag} */,
  {32'hc35375f6, 32'h41edcf7b} /* (4, 23, 28) {real, imag} */,
  {32'h4302321b, 32'hc31fda2e} /* (4, 23, 27) {real, imag} */,
  {32'h4253c9b8, 32'hc20e9856} /* (4, 23, 26) {real, imag} */,
  {32'hc20846c7, 32'h4248741c} /* (4, 23, 25) {real, imag} */,
  {32'hc271446e, 32'hc1d72cfc} /* (4, 23, 24) {real, imag} */,
  {32'h428fd996, 32'hc1803fc8} /* (4, 23, 23) {real, imag} */,
  {32'hc1da7f05, 32'h42a43c4f} /* (4, 23, 22) {real, imag} */,
  {32'h423f72cf, 32'hc2ec552a} /* (4, 23, 21) {real, imag} */,
  {32'hc1bb463f, 32'hc23e4e10} /* (4, 23, 20) {real, imag} */,
  {32'hc1afcc7e, 32'hc199d660} /* (4, 23, 19) {real, imag} */,
  {32'h4219d198, 32'hc299a902} /* (4, 23, 18) {real, imag} */,
  {32'h41d44a62, 32'h415d7646} /* (4, 23, 17) {real, imag} */,
  {32'h4211a6cf, 32'h00000000} /* (4, 23, 16) {real, imag} */,
  {32'h41d44a62, 32'hc15d7646} /* (4, 23, 15) {real, imag} */,
  {32'h4219d198, 32'h4299a902} /* (4, 23, 14) {real, imag} */,
  {32'hc1afcc7e, 32'h4199d660} /* (4, 23, 13) {real, imag} */,
  {32'hc1bb463f, 32'h423e4e10} /* (4, 23, 12) {real, imag} */,
  {32'h423f72cf, 32'h42ec552a} /* (4, 23, 11) {real, imag} */,
  {32'hc1da7f05, 32'hc2a43c4f} /* (4, 23, 10) {real, imag} */,
  {32'h428fd996, 32'h41803fc8} /* (4, 23, 9) {real, imag} */,
  {32'hc271446e, 32'h41d72cfc} /* (4, 23, 8) {real, imag} */,
  {32'hc20846c7, 32'hc248741c} /* (4, 23, 7) {real, imag} */,
  {32'h4253c9b8, 32'h420e9856} /* (4, 23, 6) {real, imag} */,
  {32'h4302321b, 32'h431fda2e} /* (4, 23, 5) {real, imag} */,
  {32'hc35375f6, 32'hc1edcf7b} /* (4, 23, 4) {real, imag} */,
  {32'hc240485c, 32'h41d9cc42} /* (4, 23, 3) {real, imag} */,
  {32'h44236956, 32'hc3493776} /* (4, 23, 2) {real, imag} */,
  {32'hc4a0d6b7, 32'h420453f8} /* (4, 23, 1) {real, imag} */,
  {32'h43160522, 32'h00000000} /* (4, 23, 0) {real, imag} */,
  {32'hc4810f06, 32'hc2c08a34} /* (4, 22, 31) {real, imag} */,
  {32'h44038c9a, 32'h43013128} /* (4, 22, 30) {real, imag} */,
  {32'hc22db437, 32'hc2b724e2} /* (4, 22, 29) {real, imag} */,
  {32'hc345778b, 32'h427e03b1} /* (4, 22, 28) {real, imag} */,
  {32'h434f2057, 32'hc1bcc592} /* (4, 22, 27) {real, imag} */,
  {32'hc1c86c02, 32'hc046d2c8} /* (4, 22, 26) {real, imag} */,
  {32'hc20b9b64, 32'hc22aa0e4} /* (4, 22, 25) {real, imag} */,
  {32'hc17b9514, 32'hc2a00803} /* (4, 22, 24) {real, imag} */,
  {32'h429cdb3d, 32'hc1a90ac6} /* (4, 22, 23) {real, imag} */,
  {32'hc1b6459a, 32'h4194b2ef} /* (4, 22, 22) {real, imag} */,
  {32'h423410e3, 32'hc3249f22} /* (4, 22, 21) {real, imag} */,
  {32'hc2348ad4, 32'hc20c745c} /* (4, 22, 20) {real, imag} */,
  {32'h42292254, 32'hc2e807ae} /* (4, 22, 19) {real, imag} */,
  {32'hc2326352, 32'hc28453ce} /* (4, 22, 18) {real, imag} */,
  {32'hc0229378, 32'h429443a2} /* (4, 22, 17) {real, imag} */,
  {32'h421d565f, 32'h00000000} /* (4, 22, 16) {real, imag} */,
  {32'hc0229378, 32'hc29443a2} /* (4, 22, 15) {real, imag} */,
  {32'hc2326352, 32'h428453ce} /* (4, 22, 14) {real, imag} */,
  {32'h42292254, 32'h42e807ae} /* (4, 22, 13) {real, imag} */,
  {32'hc2348ad4, 32'h420c745c} /* (4, 22, 12) {real, imag} */,
  {32'h423410e3, 32'h43249f22} /* (4, 22, 11) {real, imag} */,
  {32'hc1b6459a, 32'hc194b2ef} /* (4, 22, 10) {real, imag} */,
  {32'h429cdb3d, 32'h41a90ac6} /* (4, 22, 9) {real, imag} */,
  {32'hc17b9514, 32'h42a00803} /* (4, 22, 8) {real, imag} */,
  {32'hc20b9b64, 32'h422aa0e4} /* (4, 22, 7) {real, imag} */,
  {32'hc1c86c02, 32'h4046d2c8} /* (4, 22, 6) {real, imag} */,
  {32'h434f2057, 32'h41bcc592} /* (4, 22, 5) {real, imag} */,
  {32'hc345778b, 32'hc27e03b1} /* (4, 22, 4) {real, imag} */,
  {32'hc22db437, 32'h42b724e2} /* (4, 22, 3) {real, imag} */,
  {32'h44038c9a, 32'hc3013128} /* (4, 22, 2) {real, imag} */,
  {32'hc4810f06, 32'h42c08a34} /* (4, 22, 1) {real, imag} */,
  {32'h4287e7b5, 32'h00000000} /* (4, 22, 0) {real, imag} */,
  {32'hc3e42cf0, 32'hc2dd603e} /* (4, 21, 31) {real, imag} */,
  {32'h42e4abca, 32'h41a75d12} /* (4, 21, 30) {real, imag} */,
  {32'h42033b60, 32'hc25d2bdb} /* (4, 21, 29) {real, imag} */,
  {32'hc22dbad0, 32'h40e827e0} /* (4, 21, 28) {real, imag} */,
  {32'h4289c4d3, 32'hc27a191b} /* (4, 21, 27) {real, imag} */,
  {32'hc2b336bd, 32'hc2783c22} /* (4, 21, 26) {real, imag} */,
  {32'h42870a23, 32'h4235f51c} /* (4, 21, 25) {real, imag} */,
  {32'hc1bae8b9, 32'h41bc3790} /* (4, 21, 24) {real, imag} */,
  {32'h41824b9c, 32'hc27f701f} /* (4, 21, 23) {real, imag} */,
  {32'hc319c4e3, 32'hc1bed5d5} /* (4, 21, 22) {real, imag} */,
  {32'hc31a5ce0, 32'hc22942c9} /* (4, 21, 21) {real, imag} */,
  {32'h4123725c, 32'h42bdc4fa} /* (4, 21, 20) {real, imag} */,
  {32'h42d3ce5e, 32'hc180c90f} /* (4, 21, 19) {real, imag} */,
  {32'h4240fa48, 32'hc237afb5} /* (4, 21, 18) {real, imag} */,
  {32'h4247dff4, 32'hc284602a} /* (4, 21, 17) {real, imag} */,
  {32'hc2214716, 32'h00000000} /* (4, 21, 16) {real, imag} */,
  {32'h4247dff4, 32'h4284602a} /* (4, 21, 15) {real, imag} */,
  {32'h4240fa48, 32'h4237afb5} /* (4, 21, 14) {real, imag} */,
  {32'h42d3ce5e, 32'h4180c90f} /* (4, 21, 13) {real, imag} */,
  {32'h4123725c, 32'hc2bdc4fa} /* (4, 21, 12) {real, imag} */,
  {32'hc31a5ce0, 32'h422942c9} /* (4, 21, 11) {real, imag} */,
  {32'hc319c4e3, 32'h41bed5d5} /* (4, 21, 10) {real, imag} */,
  {32'h41824b9c, 32'h427f701f} /* (4, 21, 9) {real, imag} */,
  {32'hc1bae8b9, 32'hc1bc3790} /* (4, 21, 8) {real, imag} */,
  {32'h42870a23, 32'hc235f51c} /* (4, 21, 7) {real, imag} */,
  {32'hc2b336bd, 32'h42783c22} /* (4, 21, 6) {real, imag} */,
  {32'h4289c4d3, 32'h427a191b} /* (4, 21, 5) {real, imag} */,
  {32'hc22dbad0, 32'hc0e827e0} /* (4, 21, 4) {real, imag} */,
  {32'h42033b60, 32'h425d2bdb} /* (4, 21, 3) {real, imag} */,
  {32'h42e4abca, 32'hc1a75d12} /* (4, 21, 2) {real, imag} */,
  {32'hc3e42cf0, 32'h42dd603e} /* (4, 21, 1) {real, imag} */,
  {32'h43ef6b8a, 32'h00000000} /* (4, 21, 0) {real, imag} */,
  {32'h43fe0a34, 32'hc39c9f6a} /* (4, 20, 31) {real, imag} */,
  {32'hc3d4a6a2, 32'hc2a5be6a} /* (4, 20, 30) {real, imag} */,
  {32'hc212cbfe, 32'hc2bdd6c6} /* (4, 20, 29) {real, imag} */,
  {32'h42942773, 32'hc28668b2} /* (4, 20, 28) {real, imag} */,
  {32'hc3081c99, 32'hc2f25f0c} /* (4, 20, 27) {real, imag} */,
  {32'hc2230af2, 32'hc2329528} /* (4, 20, 26) {real, imag} */,
  {32'h4264f21d, 32'h431f4c9c} /* (4, 20, 25) {real, imag} */,
  {32'hc2d8a8aa, 32'hc08f8ca0} /* (4, 20, 24) {real, imag} */,
  {32'hc284b616, 32'hc23107fb} /* (4, 20, 23) {real, imag} */,
  {32'hc2d05062, 32'hc1be846c} /* (4, 20, 22) {real, imag} */,
  {32'hc2d5fe6c, 32'hc199630e} /* (4, 20, 21) {real, imag} */,
  {32'hc21790c6, 32'hc200d9b1} /* (4, 20, 20) {real, imag} */,
  {32'hc27ebfe6, 32'h428a209b} /* (4, 20, 19) {real, imag} */,
  {32'h41c3b8fc, 32'h4245dac8} /* (4, 20, 18) {real, imag} */,
  {32'h4251a810, 32'hc2a3ee98} /* (4, 20, 17) {real, imag} */,
  {32'hc21415b8, 32'h00000000} /* (4, 20, 16) {real, imag} */,
  {32'h4251a810, 32'h42a3ee98} /* (4, 20, 15) {real, imag} */,
  {32'h41c3b8fc, 32'hc245dac8} /* (4, 20, 14) {real, imag} */,
  {32'hc27ebfe6, 32'hc28a209b} /* (4, 20, 13) {real, imag} */,
  {32'hc21790c6, 32'h4200d9b1} /* (4, 20, 12) {real, imag} */,
  {32'hc2d5fe6c, 32'h4199630e} /* (4, 20, 11) {real, imag} */,
  {32'hc2d05062, 32'h41be846c} /* (4, 20, 10) {real, imag} */,
  {32'hc284b616, 32'h423107fb} /* (4, 20, 9) {real, imag} */,
  {32'hc2d8a8aa, 32'h408f8ca0} /* (4, 20, 8) {real, imag} */,
  {32'h4264f21d, 32'hc31f4c9c} /* (4, 20, 7) {real, imag} */,
  {32'hc2230af2, 32'h42329528} /* (4, 20, 6) {real, imag} */,
  {32'hc3081c99, 32'h42f25f0c} /* (4, 20, 5) {real, imag} */,
  {32'h42942773, 32'h428668b2} /* (4, 20, 4) {real, imag} */,
  {32'hc212cbfe, 32'h42bdd6c6} /* (4, 20, 3) {real, imag} */,
  {32'hc3d4a6a2, 32'h42a5be6a} /* (4, 20, 2) {real, imag} */,
  {32'h43fe0a34, 32'h439c9f6a} /* (4, 20, 1) {real, imag} */,
  {32'h448a0758, 32'h00000000} /* (4, 20, 0) {real, imag} */,
  {32'h4451b273, 32'hc32fb1b4} /* (4, 19, 31) {real, imag} */,
  {32'hc40d3c5f, 32'h417b44e8} /* (4, 19, 30) {real, imag} */,
  {32'hc297ad2a, 32'hc16155e6} /* (4, 19, 29) {real, imag} */,
  {32'h4230f0a0, 32'hc3298242} /* (4, 19, 28) {real, imag} */,
  {32'hc2deee80, 32'hc20eb7d0} /* (4, 19, 27) {real, imag} */,
  {32'hc2022b06, 32'hc2c7e0b0} /* (4, 19, 26) {real, imag} */,
  {32'h42602714, 32'h3da33800} /* (4, 19, 25) {real, imag} */,
  {32'hc10a9d2c, 32'h419aa724} /* (4, 19, 24) {real, imag} */,
  {32'h4281477b, 32'h4112d9c6} /* (4, 19, 23) {real, imag} */,
  {32'h42004a48, 32'hc10e65e0} /* (4, 19, 22) {real, imag} */,
  {32'hc2675cb8, 32'h42dd0b4d} /* (4, 19, 21) {real, imag} */,
  {32'h41817fa4, 32'h40eaa6b0} /* (4, 19, 20) {real, imag} */,
  {32'h409dd17c, 32'h42990436} /* (4, 19, 19) {real, imag} */,
  {32'h42ab7870, 32'h4289e9f6} /* (4, 19, 18) {real, imag} */,
  {32'hc1ca6c8a, 32'h42ae2fc5} /* (4, 19, 17) {real, imag} */,
  {32'h429a3dcd, 32'h00000000} /* (4, 19, 16) {real, imag} */,
  {32'hc1ca6c8a, 32'hc2ae2fc5} /* (4, 19, 15) {real, imag} */,
  {32'h42ab7870, 32'hc289e9f6} /* (4, 19, 14) {real, imag} */,
  {32'h409dd17c, 32'hc2990436} /* (4, 19, 13) {real, imag} */,
  {32'h41817fa4, 32'hc0eaa6b0} /* (4, 19, 12) {real, imag} */,
  {32'hc2675cb8, 32'hc2dd0b4d} /* (4, 19, 11) {real, imag} */,
  {32'h42004a48, 32'h410e65e0} /* (4, 19, 10) {real, imag} */,
  {32'h4281477b, 32'hc112d9c6} /* (4, 19, 9) {real, imag} */,
  {32'hc10a9d2c, 32'hc19aa724} /* (4, 19, 8) {real, imag} */,
  {32'h42602714, 32'hbda33800} /* (4, 19, 7) {real, imag} */,
  {32'hc2022b06, 32'h42c7e0b0} /* (4, 19, 6) {real, imag} */,
  {32'hc2deee80, 32'h420eb7d0} /* (4, 19, 5) {real, imag} */,
  {32'h4230f0a0, 32'h43298242} /* (4, 19, 4) {real, imag} */,
  {32'hc297ad2a, 32'h416155e6} /* (4, 19, 3) {real, imag} */,
  {32'hc40d3c5f, 32'hc17b44e8} /* (4, 19, 2) {real, imag} */,
  {32'h4451b273, 32'h432fb1b4} /* (4, 19, 1) {real, imag} */,
  {32'h44563718, 32'h00000000} /* (4, 19, 0) {real, imag} */,
  {32'h446056fc, 32'hc2e8e2c8} /* (4, 18, 31) {real, imag} */,
  {32'hc408b655, 32'h435f29c7} /* (4, 18, 30) {real, imag} */,
  {32'hc2b1adb1, 32'hc2b44668} /* (4, 18, 29) {real, imag} */,
  {32'h42b09169, 32'hc31bdc24} /* (4, 18, 28) {real, imag} */,
  {32'hc31911f4, 32'hc2205754} /* (4, 18, 27) {real, imag} */,
  {32'h4200455c, 32'hbfb82700} /* (4, 18, 26) {real, imag} */,
  {32'h427e2b9c, 32'hc17af444} /* (4, 18, 25) {real, imag} */,
  {32'hc1ed06f6, 32'h43009c72} /* (4, 18, 24) {real, imag} */,
  {32'hc0937ed0, 32'hc059cb98} /* (4, 18, 23) {real, imag} */,
  {32'hc2646a1a, 32'hc2814d42} /* (4, 18, 22) {real, imag} */,
  {32'h4161ded8, 32'h43032cce} /* (4, 18, 21) {real, imag} */,
  {32'hc24fc546, 32'h41ade3fa} /* (4, 18, 20) {real, imag} */,
  {32'hc2749f61, 32'hc1de2356} /* (4, 18, 19) {real, imag} */,
  {32'h4222f122, 32'h42096e1e} /* (4, 18, 18) {real, imag} */,
  {32'hc19b4a9e, 32'hc2387abb} /* (4, 18, 17) {real, imag} */,
  {32'h42433779, 32'h00000000} /* (4, 18, 16) {real, imag} */,
  {32'hc19b4a9e, 32'h42387abb} /* (4, 18, 15) {real, imag} */,
  {32'h4222f122, 32'hc2096e1e} /* (4, 18, 14) {real, imag} */,
  {32'hc2749f61, 32'h41de2356} /* (4, 18, 13) {real, imag} */,
  {32'hc24fc546, 32'hc1ade3fa} /* (4, 18, 12) {real, imag} */,
  {32'h4161ded8, 32'hc3032cce} /* (4, 18, 11) {real, imag} */,
  {32'hc2646a1a, 32'h42814d42} /* (4, 18, 10) {real, imag} */,
  {32'hc0937ed0, 32'h4059cb98} /* (4, 18, 9) {real, imag} */,
  {32'hc1ed06f6, 32'hc3009c72} /* (4, 18, 8) {real, imag} */,
  {32'h427e2b9c, 32'h417af444} /* (4, 18, 7) {real, imag} */,
  {32'h4200455c, 32'h3fb82700} /* (4, 18, 6) {real, imag} */,
  {32'hc31911f4, 32'h42205754} /* (4, 18, 5) {real, imag} */,
  {32'h42b09169, 32'h431bdc24} /* (4, 18, 4) {real, imag} */,
  {32'hc2b1adb1, 32'h42b44668} /* (4, 18, 3) {real, imag} */,
  {32'hc408b655, 32'hc35f29c7} /* (4, 18, 2) {real, imag} */,
  {32'h446056fc, 32'h42e8e2c8} /* (4, 18, 1) {real, imag} */,
  {32'h445664eb, 32'h00000000} /* (4, 18, 0) {real, imag} */,
  {32'h4480949d, 32'hc2b42c08} /* (4, 17, 31) {real, imag} */,
  {32'hc41023fa, 32'h436842d1} /* (4, 17, 30) {real, imag} */,
  {32'hc2bb9ae4, 32'h40047aa0} /* (4, 17, 29) {real, imag} */,
  {32'h41320538, 32'hc26793ac} /* (4, 17, 28) {real, imag} */,
  {32'hc3304680, 32'hc043a980} /* (4, 17, 27) {real, imag} */,
  {32'hc02bf558, 32'hc20cdb24} /* (4, 17, 26) {real, imag} */,
  {32'h42e63e9a, 32'hc27e87ee} /* (4, 17, 25) {real, imag} */,
  {32'hc32a3d83, 32'h42c8e8b8} /* (4, 17, 24) {real, imag} */,
  {32'hc241ce10, 32'hc205dace} /* (4, 17, 23) {real, imag} */,
  {32'hc274b834, 32'h41c0dc08} /* (4, 17, 22) {real, imag} */,
  {32'hc1e0a273, 32'h4202b2dd} /* (4, 17, 21) {real, imag} */,
  {32'hc1dd34c6, 32'hc2b36450} /* (4, 17, 20) {real, imag} */,
  {32'h423823e4, 32'h41b935ad} /* (4, 17, 19) {real, imag} */,
  {32'h3f2e22e0, 32'h42b8e817} /* (4, 17, 18) {real, imag} */,
  {32'hc264f0a0, 32'h403a0240} /* (4, 17, 17) {real, imag} */,
  {32'h416ae786, 32'h00000000} /* (4, 17, 16) {real, imag} */,
  {32'hc264f0a0, 32'hc03a0240} /* (4, 17, 15) {real, imag} */,
  {32'h3f2e22e0, 32'hc2b8e817} /* (4, 17, 14) {real, imag} */,
  {32'h423823e4, 32'hc1b935ad} /* (4, 17, 13) {real, imag} */,
  {32'hc1dd34c6, 32'h42b36450} /* (4, 17, 12) {real, imag} */,
  {32'hc1e0a273, 32'hc202b2dd} /* (4, 17, 11) {real, imag} */,
  {32'hc274b834, 32'hc1c0dc08} /* (4, 17, 10) {real, imag} */,
  {32'hc241ce10, 32'h4205dace} /* (4, 17, 9) {real, imag} */,
  {32'hc32a3d83, 32'hc2c8e8b8} /* (4, 17, 8) {real, imag} */,
  {32'h42e63e9a, 32'h427e87ee} /* (4, 17, 7) {real, imag} */,
  {32'hc02bf558, 32'h420cdb24} /* (4, 17, 6) {real, imag} */,
  {32'hc3304680, 32'h4043a980} /* (4, 17, 5) {real, imag} */,
  {32'h41320538, 32'h426793ac} /* (4, 17, 4) {real, imag} */,
  {32'hc2bb9ae4, 32'hc0047aa0} /* (4, 17, 3) {real, imag} */,
  {32'hc41023fa, 32'hc36842d1} /* (4, 17, 2) {real, imag} */,
  {32'h4480949d, 32'h42b42c08} /* (4, 17, 1) {real, imag} */,
  {32'h444c2e3f, 32'h00000000} /* (4, 17, 0) {real, imag} */,
  {32'h4483c284, 32'hc3576417} /* (4, 16, 31) {real, imag} */,
  {32'hc41ea174, 32'h434d3afc} /* (4, 16, 30) {real, imag} */,
  {32'hc19f5451, 32'hc08539b0} /* (4, 16, 29) {real, imag} */,
  {32'h43081b22, 32'hc2f07758} /* (4, 16, 28) {real, imag} */,
  {32'hc2a640fc, 32'h43205a7c} /* (4, 16, 27) {real, imag} */,
  {32'hc2232c34, 32'hc1e6898b} /* (4, 16, 26) {real, imag} */,
  {32'h41b84d3a, 32'hc30a104e} /* (4, 16, 25) {real, imag} */,
  {32'hc2b5f66c, 32'h42f4851f} /* (4, 16, 24) {real, imag} */,
  {32'h4266a1ad, 32'hc12be414} /* (4, 16, 23) {real, imag} */,
  {32'h41925283, 32'h42a6bb10} /* (4, 16, 22) {real, imag} */,
  {32'h42258732, 32'hc245a170} /* (4, 16, 21) {real, imag} */,
  {32'h42247930, 32'hc270af54} /* (4, 16, 20) {real, imag} */,
  {32'h426f8f8c, 32'hc1984ee6} /* (4, 16, 19) {real, imag} */,
  {32'h423eb334, 32'h40be6564} /* (4, 16, 18) {real, imag} */,
  {32'hc15c44c1, 32'hc22b5a75} /* (4, 16, 17) {real, imag} */,
  {32'hc1db9c98, 32'h00000000} /* (4, 16, 16) {real, imag} */,
  {32'hc15c44c1, 32'h422b5a75} /* (4, 16, 15) {real, imag} */,
  {32'h423eb334, 32'hc0be6564} /* (4, 16, 14) {real, imag} */,
  {32'h426f8f8c, 32'h41984ee6} /* (4, 16, 13) {real, imag} */,
  {32'h42247930, 32'h4270af54} /* (4, 16, 12) {real, imag} */,
  {32'h42258732, 32'h4245a170} /* (4, 16, 11) {real, imag} */,
  {32'h41925283, 32'hc2a6bb10} /* (4, 16, 10) {real, imag} */,
  {32'h4266a1ad, 32'h412be414} /* (4, 16, 9) {real, imag} */,
  {32'hc2b5f66c, 32'hc2f4851f} /* (4, 16, 8) {real, imag} */,
  {32'h41b84d3a, 32'h430a104e} /* (4, 16, 7) {real, imag} */,
  {32'hc2232c34, 32'h41e6898b} /* (4, 16, 6) {real, imag} */,
  {32'hc2a640fc, 32'hc3205a7c} /* (4, 16, 5) {real, imag} */,
  {32'h43081b22, 32'h42f07758} /* (4, 16, 4) {real, imag} */,
  {32'hc19f5451, 32'h408539b0} /* (4, 16, 3) {real, imag} */,
  {32'hc41ea174, 32'hc34d3afc} /* (4, 16, 2) {real, imag} */,
  {32'h4483c284, 32'h43576417} /* (4, 16, 1) {real, imag} */,
  {32'h442344fe, 32'h00000000} /* (4, 16, 0) {real, imag} */,
  {32'h447f9516, 32'hc3cee3e4} /* (4, 15, 31) {real, imag} */,
  {32'hc417e74a, 32'h42a12162} /* (4, 15, 30) {real, imag} */,
  {32'h42c58430, 32'hc3065016} /* (4, 15, 29) {real, imag} */,
  {32'h434ddcec, 32'hc251f126} /* (4, 15, 28) {real, imag} */,
  {32'hc38b6c10, 32'h4301b739} /* (4, 15, 27) {real, imag} */,
  {32'h4227467a, 32'h42646a08} /* (4, 15, 26) {real, imag} */,
  {32'h41eab590, 32'h410bfb2e} /* (4, 15, 25) {real, imag} */,
  {32'hc2670dfc, 32'h42490f99} /* (4, 15, 24) {real, imag} */,
  {32'h4238d08c, 32'h42ad368a} /* (4, 15, 23) {real, imag} */,
  {32'h41a1c524, 32'h421fe158} /* (4, 15, 22) {real, imag} */,
  {32'h3ff6aff0, 32'h425b812d} /* (4, 15, 21) {real, imag} */,
  {32'h40f26288, 32'h42816acc} /* (4, 15, 20) {real, imag} */,
  {32'hc140d5a6, 32'h40ef33a4} /* (4, 15, 19) {real, imag} */,
  {32'h425de5cc, 32'h42b84365} /* (4, 15, 18) {real, imag} */,
  {32'h3e55d080, 32'hc2c031b9} /* (4, 15, 17) {real, imag} */,
  {32'h42541b7e, 32'h00000000} /* (4, 15, 16) {real, imag} */,
  {32'h3e55d080, 32'h42c031b9} /* (4, 15, 15) {real, imag} */,
  {32'h425de5cc, 32'hc2b84365} /* (4, 15, 14) {real, imag} */,
  {32'hc140d5a6, 32'hc0ef33a4} /* (4, 15, 13) {real, imag} */,
  {32'h40f26288, 32'hc2816acc} /* (4, 15, 12) {real, imag} */,
  {32'h3ff6aff0, 32'hc25b812d} /* (4, 15, 11) {real, imag} */,
  {32'h41a1c524, 32'hc21fe158} /* (4, 15, 10) {real, imag} */,
  {32'h4238d08c, 32'hc2ad368a} /* (4, 15, 9) {real, imag} */,
  {32'hc2670dfc, 32'hc2490f99} /* (4, 15, 8) {real, imag} */,
  {32'h41eab590, 32'hc10bfb2e} /* (4, 15, 7) {real, imag} */,
  {32'h4227467a, 32'hc2646a08} /* (4, 15, 6) {real, imag} */,
  {32'hc38b6c10, 32'hc301b739} /* (4, 15, 5) {real, imag} */,
  {32'h434ddcec, 32'h4251f126} /* (4, 15, 4) {real, imag} */,
  {32'h42c58430, 32'h43065016} /* (4, 15, 3) {real, imag} */,
  {32'hc417e74a, 32'hc2a12162} /* (4, 15, 2) {real, imag} */,
  {32'h447f9516, 32'h43cee3e4} /* (4, 15, 1) {real, imag} */,
  {32'h442a43e5, 32'h00000000} /* (4, 15, 0) {real, imag} */,
  {32'h44808084, 32'hc38715ac} /* (4, 14, 31) {real, imag} */,
  {32'hc40cbedf, 32'hc1a1ba48} /* (4, 14, 30) {real, imag} */,
  {32'h42f6e325, 32'hc3523594} /* (4, 14, 29) {real, imag} */,
  {32'h42e313ab, 32'hc2ee9fdf} /* (4, 14, 28) {real, imag} */,
  {32'hc286aa61, 32'h4305b187} /* (4, 14, 27) {real, imag} */,
  {32'h42a34e74, 32'h42bd3420} /* (4, 14, 26) {real, imag} */,
  {32'h42c51ae2, 32'hc12a49ec} /* (4, 14, 25) {real, imag} */,
  {32'hc1296a4d, 32'h41cbdf5c} /* (4, 14, 24) {real, imag} */,
  {32'h429237bb, 32'h421a3ed6} /* (4, 14, 23) {real, imag} */,
  {32'h422c3874, 32'hc1873a5e} /* (4, 14, 22) {real, imag} */,
  {32'hc30c2d8e, 32'h4179663c} /* (4, 14, 21) {real, imag} */,
  {32'hc23c1714, 32'h41923054} /* (4, 14, 20) {real, imag} */,
  {32'hc2d0bace, 32'hbfdc05c0} /* (4, 14, 19) {real, imag} */,
  {32'h40b0409c, 32'h42647810} /* (4, 14, 18) {real, imag} */,
  {32'hc2b30ca0, 32'h424f187d} /* (4, 14, 17) {real, imag} */,
  {32'hc22c5a5f, 32'h00000000} /* (4, 14, 16) {real, imag} */,
  {32'hc2b30ca0, 32'hc24f187d} /* (4, 14, 15) {real, imag} */,
  {32'h40b0409c, 32'hc2647810} /* (4, 14, 14) {real, imag} */,
  {32'hc2d0bace, 32'h3fdc05c0} /* (4, 14, 13) {real, imag} */,
  {32'hc23c1714, 32'hc1923054} /* (4, 14, 12) {real, imag} */,
  {32'hc30c2d8e, 32'hc179663c} /* (4, 14, 11) {real, imag} */,
  {32'h422c3874, 32'h41873a5e} /* (4, 14, 10) {real, imag} */,
  {32'h429237bb, 32'hc21a3ed6} /* (4, 14, 9) {real, imag} */,
  {32'hc1296a4d, 32'hc1cbdf5c} /* (4, 14, 8) {real, imag} */,
  {32'h42c51ae2, 32'h412a49ec} /* (4, 14, 7) {real, imag} */,
  {32'h42a34e74, 32'hc2bd3420} /* (4, 14, 6) {real, imag} */,
  {32'hc286aa61, 32'hc305b187} /* (4, 14, 5) {real, imag} */,
  {32'h42e313ab, 32'h42ee9fdf} /* (4, 14, 4) {real, imag} */,
  {32'h42f6e325, 32'h43523594} /* (4, 14, 3) {real, imag} */,
  {32'hc40cbedf, 32'h41a1ba48} /* (4, 14, 2) {real, imag} */,
  {32'h44808084, 32'h438715ac} /* (4, 14, 1) {real, imag} */,
  {32'h4434b3a1, 32'h00000000} /* (4, 14, 0) {real, imag} */,
  {32'h4483c8b6, 32'hc37c5a98} /* (4, 13, 31) {real, imag} */,
  {32'hc3dff9f6, 32'hc28dd99d} /* (4, 13, 30) {real, imag} */,
  {32'h4324f51c, 32'h4237fd1a} /* (4, 13, 29) {real, imag} */,
  {32'h42c9ff3a, 32'hc291b028} /* (4, 13, 28) {real, imag} */,
  {32'hc2ec4474, 32'h437e86e4} /* (4, 13, 27) {real, imag} */,
  {32'h43490994, 32'h42bf517c} /* (4, 13, 26) {real, imag} */,
  {32'hc0a9a4fc, 32'hc1ae6c6f} /* (4, 13, 25) {real, imag} */,
  {32'hc2ae2e22, 32'h4216785a} /* (4, 13, 24) {real, imag} */,
  {32'h427658d4, 32'h413c7b22} /* (4, 13, 23) {real, imag} */,
  {32'hc1dd2a3d, 32'hc2803444} /* (4, 13, 22) {real, imag} */,
  {32'h41a20cf0, 32'h42e4c13b} /* (4, 13, 21) {real, imag} */,
  {32'h429cbe62, 32'hc2725ff2} /* (4, 13, 20) {real, imag} */,
  {32'h41c81197, 32'hc2593cd3} /* (4, 13, 19) {real, imag} */,
  {32'h41f2a07c, 32'h4111364e} /* (4, 13, 18) {real, imag} */,
  {32'hc0cfee8e, 32'hc1d0e23c} /* (4, 13, 17) {real, imag} */,
  {32'h4222c33a, 32'h00000000} /* (4, 13, 16) {real, imag} */,
  {32'hc0cfee8e, 32'h41d0e23c} /* (4, 13, 15) {real, imag} */,
  {32'h41f2a07c, 32'hc111364e} /* (4, 13, 14) {real, imag} */,
  {32'h41c81197, 32'h42593cd3} /* (4, 13, 13) {real, imag} */,
  {32'h429cbe62, 32'h42725ff2} /* (4, 13, 12) {real, imag} */,
  {32'h41a20cf0, 32'hc2e4c13b} /* (4, 13, 11) {real, imag} */,
  {32'hc1dd2a3d, 32'h42803444} /* (4, 13, 10) {real, imag} */,
  {32'h427658d4, 32'hc13c7b22} /* (4, 13, 9) {real, imag} */,
  {32'hc2ae2e22, 32'hc216785a} /* (4, 13, 8) {real, imag} */,
  {32'hc0a9a4fc, 32'h41ae6c6f} /* (4, 13, 7) {real, imag} */,
  {32'h43490994, 32'hc2bf517c} /* (4, 13, 6) {real, imag} */,
  {32'hc2ec4474, 32'hc37e86e4} /* (4, 13, 5) {real, imag} */,
  {32'h42c9ff3a, 32'h4291b028} /* (4, 13, 4) {real, imag} */,
  {32'h4324f51c, 32'hc237fd1a} /* (4, 13, 3) {real, imag} */,
  {32'hc3dff9f6, 32'h428dd99d} /* (4, 13, 2) {real, imag} */,
  {32'h4483c8b6, 32'h437c5a98} /* (4, 13, 1) {real, imag} */,
  {32'h441dd89a, 32'h00000000} /* (4, 13, 0) {real, imag} */,
  {32'h44626e9e, 32'hc3629d19} /* (4, 12, 31) {real, imag} */,
  {32'hc3e1ef8a, 32'hc20a021b} /* (4, 12, 30) {real, imag} */,
  {32'h43297e28, 32'h42aac09c} /* (4, 12, 29) {real, imag} */,
  {32'h42a3cf69, 32'hc27b949c} /* (4, 12, 28) {real, imag} */,
  {32'hc37601f9, 32'h42a79694} /* (4, 12, 27) {real, imag} */,
  {32'h42bc5f19, 32'h42b7f0ce} /* (4, 12, 26) {real, imag} */,
  {32'h41beabb6, 32'h41e3c684} /* (4, 12, 25) {real, imag} */,
  {32'hc27ca46d, 32'h4286356c} /* (4, 12, 24) {real, imag} */,
  {32'h4286e81a, 32'hbd511000} /* (4, 12, 23) {real, imag} */,
  {32'h402fbcb0, 32'h41793bc4} /* (4, 12, 22) {real, imag} */,
  {32'hc1f71938, 32'h42d80e8a} /* (4, 12, 21) {real, imag} */,
  {32'h400584b8, 32'hc225280b} /* (4, 12, 20) {real, imag} */,
  {32'h41abe06b, 32'hc22b9f62} /* (4, 12, 19) {real, imag} */,
  {32'h412ead40, 32'hc2852ab8} /* (4, 12, 18) {real, imag} */,
  {32'h410371ea, 32'h41c69922} /* (4, 12, 17) {real, imag} */,
  {32'h42ded54c, 32'h00000000} /* (4, 12, 16) {real, imag} */,
  {32'h410371ea, 32'hc1c69922} /* (4, 12, 15) {real, imag} */,
  {32'h412ead40, 32'h42852ab8} /* (4, 12, 14) {real, imag} */,
  {32'h41abe06b, 32'h422b9f62} /* (4, 12, 13) {real, imag} */,
  {32'h400584b8, 32'h4225280b} /* (4, 12, 12) {real, imag} */,
  {32'hc1f71938, 32'hc2d80e8a} /* (4, 12, 11) {real, imag} */,
  {32'h402fbcb0, 32'hc1793bc4} /* (4, 12, 10) {real, imag} */,
  {32'h4286e81a, 32'h3d511000} /* (4, 12, 9) {real, imag} */,
  {32'hc27ca46d, 32'hc286356c} /* (4, 12, 8) {real, imag} */,
  {32'h41beabb6, 32'hc1e3c684} /* (4, 12, 7) {real, imag} */,
  {32'h42bc5f19, 32'hc2b7f0ce} /* (4, 12, 6) {real, imag} */,
  {32'hc37601f9, 32'hc2a79694} /* (4, 12, 5) {real, imag} */,
  {32'h42a3cf69, 32'h427b949c} /* (4, 12, 4) {real, imag} */,
  {32'h43297e28, 32'hc2aac09c} /* (4, 12, 3) {real, imag} */,
  {32'hc3e1ef8a, 32'h420a021b} /* (4, 12, 2) {real, imag} */,
  {32'h44626e9e, 32'h43629d19} /* (4, 12, 1) {real, imag} */,
  {32'h44335a46, 32'h00000000} /* (4, 12, 0) {real, imag} */,
  {32'h443380d2, 32'hc362c373} /* (4, 11, 31) {real, imag} */,
  {32'hc3b58202, 32'hc1ae7276} /* (4, 11, 30) {real, imag} */,
  {32'h4323f03d, 32'hc1c1df66} /* (4, 11, 29) {real, imag} */,
  {32'h42447898, 32'hc231b898} /* (4, 11, 28) {real, imag} */,
  {32'hc350f924, 32'h42a33230} /* (4, 11, 27) {real, imag} */,
  {32'h4332660a, 32'h425fe128} /* (4, 11, 26) {real, imag} */,
  {32'h422a5b9a, 32'h4274f5e8} /* (4, 11, 25) {real, imag} */,
  {32'hc23a7174, 32'h41fb1908} /* (4, 11, 24) {real, imag} */,
  {32'hc22db3ba, 32'hc219b641} /* (4, 11, 23) {real, imag} */,
  {32'h4301169f, 32'h41d33d6b} /* (4, 11, 22) {real, imag} */,
  {32'hc29241ad, 32'h41e77fbe} /* (4, 11, 21) {real, imag} */,
  {32'hc2344435, 32'h40df90a0} /* (4, 11, 20) {real, imag} */,
  {32'h4162efcc, 32'h427585ce} /* (4, 11, 19) {real, imag} */,
  {32'h40f094a4, 32'h42f11a9a} /* (4, 11, 18) {real, imag} */,
  {32'hc1dfb640, 32'hc143d8a2} /* (4, 11, 17) {real, imag} */,
  {32'h420379b0, 32'h00000000} /* (4, 11, 16) {real, imag} */,
  {32'hc1dfb640, 32'h4143d8a2} /* (4, 11, 15) {real, imag} */,
  {32'h40f094a4, 32'hc2f11a9a} /* (4, 11, 14) {real, imag} */,
  {32'h4162efcc, 32'hc27585ce} /* (4, 11, 13) {real, imag} */,
  {32'hc2344435, 32'hc0df90a0} /* (4, 11, 12) {real, imag} */,
  {32'hc29241ad, 32'hc1e77fbe} /* (4, 11, 11) {real, imag} */,
  {32'h4301169f, 32'hc1d33d6b} /* (4, 11, 10) {real, imag} */,
  {32'hc22db3ba, 32'h4219b641} /* (4, 11, 9) {real, imag} */,
  {32'hc23a7174, 32'hc1fb1908} /* (4, 11, 8) {real, imag} */,
  {32'h422a5b9a, 32'hc274f5e8} /* (4, 11, 7) {real, imag} */,
  {32'h4332660a, 32'hc25fe128} /* (4, 11, 6) {real, imag} */,
  {32'hc350f924, 32'hc2a33230} /* (4, 11, 5) {real, imag} */,
  {32'h42447898, 32'h4231b898} /* (4, 11, 4) {real, imag} */,
  {32'h4323f03d, 32'h41c1df66} /* (4, 11, 3) {real, imag} */,
  {32'hc3b58202, 32'h41ae7276} /* (4, 11, 2) {real, imag} */,
  {32'h443380d2, 32'h4362c373} /* (4, 11, 1) {real, imag} */,
  {32'h441a2f81, 32'h00000000} /* (4, 11, 0) {real, imag} */,
  {32'hc2c5ce50, 32'hc301ce7f} /* (4, 10, 31) {real, imag} */,
  {32'h435598de, 32'hc2b753a7} /* (4, 10, 30) {real, imag} */,
  {32'h43169152, 32'hc1863946} /* (4, 10, 29) {real, imag} */,
  {32'hc28e3d8a, 32'hc1d54892} /* (4, 10, 28) {real, imag} */,
  {32'h42466534, 32'hc2b59702} /* (4, 10, 27) {real, imag} */,
  {32'h42ea221c, 32'hc209f3d8} /* (4, 10, 26) {real, imag} */,
  {32'hc2eb29b4, 32'h42fbbc20} /* (4, 10, 25) {real, imag} */,
  {32'h424ca7c9, 32'hc24615a6} /* (4, 10, 24) {real, imag} */,
  {32'hc2cdf8f5, 32'h42bdf1d4} /* (4, 10, 23) {real, imag} */,
  {32'hc0a5e1e6, 32'hc1bb63ed} /* (4, 10, 22) {real, imag} */,
  {32'hc1f94b2b, 32'hc29f7a5d} /* (4, 10, 21) {real, imag} */,
  {32'h41f8bb98, 32'h42ccfe5a} /* (4, 10, 20) {real, imag} */,
  {32'hc0e5a9b8, 32'hc25a66d5} /* (4, 10, 19) {real, imag} */,
  {32'hc299f92f, 32'h40e89978} /* (4, 10, 18) {real, imag} */,
  {32'h4208f0d8, 32'h424e09d0} /* (4, 10, 17) {real, imag} */,
  {32'hc19861fe, 32'h00000000} /* (4, 10, 16) {real, imag} */,
  {32'h4208f0d8, 32'hc24e09d0} /* (4, 10, 15) {real, imag} */,
  {32'hc299f92f, 32'hc0e89978} /* (4, 10, 14) {real, imag} */,
  {32'hc0e5a9b8, 32'h425a66d5} /* (4, 10, 13) {real, imag} */,
  {32'h41f8bb98, 32'hc2ccfe5a} /* (4, 10, 12) {real, imag} */,
  {32'hc1f94b2b, 32'h429f7a5d} /* (4, 10, 11) {real, imag} */,
  {32'hc0a5e1e6, 32'h41bb63ed} /* (4, 10, 10) {real, imag} */,
  {32'hc2cdf8f5, 32'hc2bdf1d4} /* (4, 10, 9) {real, imag} */,
  {32'h424ca7c9, 32'h424615a6} /* (4, 10, 8) {real, imag} */,
  {32'hc2eb29b4, 32'hc2fbbc20} /* (4, 10, 7) {real, imag} */,
  {32'h42ea221c, 32'h4209f3d8} /* (4, 10, 6) {real, imag} */,
  {32'h42466534, 32'h42b59702} /* (4, 10, 5) {real, imag} */,
  {32'hc28e3d8a, 32'h41d54892} /* (4, 10, 4) {real, imag} */,
  {32'h43169152, 32'h41863946} /* (4, 10, 3) {real, imag} */,
  {32'h435598de, 32'h42b753a7} /* (4, 10, 2) {real, imag} */,
  {32'hc2c5ce50, 32'h4301ce7f} /* (4, 10, 1) {real, imag} */,
  {32'hc25b9da2, 32'h00000000} /* (4, 10, 0) {real, imag} */,
  {32'hc41daf98, 32'hc2a39b8e} /* (4, 9, 31) {real, imag} */,
  {32'h43dd0fd5, 32'hc0901ff0} /* (4, 9, 30) {real, imag} */,
  {32'h42a36cc4, 32'hc21286e9} /* (4, 9, 29) {real, imag} */,
  {32'hc2dd836f, 32'h422a0302} /* (4, 9, 28) {real, imag} */,
  {32'h434c6487, 32'hc3294f4e} /* (4, 9, 27) {real, imag} */,
  {32'h42e97880, 32'hc208d3b4} /* (4, 9, 26) {real, imag} */,
  {32'hc283c132, 32'h424de248} /* (4, 9, 25) {real, imag} */,
  {32'h426858bc, 32'hc2b31c6e} /* (4, 9, 24) {real, imag} */,
  {32'h42013860, 32'h415ed4b8} /* (4, 9, 23) {real, imag} */,
  {32'h4187e13d, 32'h41e0d6e4} /* (4, 9, 22) {real, imag} */,
  {32'hbe001f00, 32'hc14f6140} /* (4, 9, 21) {real, imag} */,
  {32'hc1c67e53, 32'h429bfc1d} /* (4, 9, 20) {real, imag} */,
  {32'h4218058f, 32'h4294eab8} /* (4, 9, 19) {real, imag} */,
  {32'hc2629840, 32'hc25c6d4f} /* (4, 9, 18) {real, imag} */,
  {32'hc2c54ed2, 32'h421e5b8e} /* (4, 9, 17) {real, imag} */,
  {32'h4289d0fa, 32'h00000000} /* (4, 9, 16) {real, imag} */,
  {32'hc2c54ed2, 32'hc21e5b8e} /* (4, 9, 15) {real, imag} */,
  {32'hc2629840, 32'h425c6d4f} /* (4, 9, 14) {real, imag} */,
  {32'h4218058f, 32'hc294eab8} /* (4, 9, 13) {real, imag} */,
  {32'hc1c67e53, 32'hc29bfc1d} /* (4, 9, 12) {real, imag} */,
  {32'hbe001f00, 32'h414f6140} /* (4, 9, 11) {real, imag} */,
  {32'h4187e13d, 32'hc1e0d6e4} /* (4, 9, 10) {real, imag} */,
  {32'h42013860, 32'hc15ed4b8} /* (4, 9, 9) {real, imag} */,
  {32'h426858bc, 32'h42b31c6e} /* (4, 9, 8) {real, imag} */,
  {32'hc283c132, 32'hc24de248} /* (4, 9, 7) {real, imag} */,
  {32'h42e97880, 32'h4208d3b4} /* (4, 9, 6) {real, imag} */,
  {32'h434c6487, 32'h43294f4e} /* (4, 9, 5) {real, imag} */,
  {32'hc2dd836f, 32'hc22a0302} /* (4, 9, 4) {real, imag} */,
  {32'h42a36cc4, 32'h421286e9} /* (4, 9, 3) {real, imag} */,
  {32'h43dd0fd5, 32'h40901ff0} /* (4, 9, 2) {real, imag} */,
  {32'hc41daf98, 32'h42a39b8e} /* (4, 9, 1) {real, imag} */,
  {32'hc2f1793c, 32'h00000000} /* (4, 9, 0) {real, imag} */,
  {32'hc44c0b48, 32'hc2ddaa3a} /* (4, 8, 31) {real, imag} */,
  {32'h440843b4, 32'h42bafe97} /* (4, 8, 30) {real, imag} */,
  {32'h43181eb1, 32'hc294ea3a} /* (4, 8, 29) {real, imag} */,
  {32'h409028c0, 32'h410a057e} /* (4, 8, 28) {real, imag} */,
  {32'h42e5fea1, 32'hc2ebd2ff} /* (4, 8, 27) {real, imag} */,
  {32'h420d9c72, 32'h42797924} /* (4, 8, 26) {real, imag} */,
  {32'hc2d4fa74, 32'h420e8730} /* (4, 8, 25) {real, imag} */,
  {32'h423d286e, 32'hc30e981a} /* (4, 8, 24) {real, imag} */,
  {32'hc24246f3, 32'hc1599cc4} /* (4, 8, 23) {real, imag} */,
  {32'h3efdb700, 32'hc296cc38} /* (4, 8, 22) {real, imag} */,
  {32'h421a7542, 32'h42c15ff5} /* (4, 8, 21) {real, imag} */,
  {32'hc2806722, 32'hc2abf0a2} /* (4, 8, 20) {real, imag} */,
  {32'h4292bcef, 32'hc18edf48} /* (4, 8, 19) {real, imag} */,
  {32'h4210208c, 32'h3ff615c0} /* (4, 8, 18) {real, imag} */,
  {32'hc03d8934, 32'h418f6b7b} /* (4, 8, 17) {real, imag} */,
  {32'hc1e29906, 32'h00000000} /* (4, 8, 16) {real, imag} */,
  {32'hc03d8934, 32'hc18f6b7b} /* (4, 8, 15) {real, imag} */,
  {32'h4210208c, 32'hbff615c0} /* (4, 8, 14) {real, imag} */,
  {32'h4292bcef, 32'h418edf48} /* (4, 8, 13) {real, imag} */,
  {32'hc2806722, 32'h42abf0a2} /* (4, 8, 12) {real, imag} */,
  {32'h421a7542, 32'hc2c15ff5} /* (4, 8, 11) {real, imag} */,
  {32'h3efdb700, 32'h4296cc38} /* (4, 8, 10) {real, imag} */,
  {32'hc24246f3, 32'h41599cc4} /* (4, 8, 9) {real, imag} */,
  {32'h423d286e, 32'h430e981a} /* (4, 8, 8) {real, imag} */,
  {32'hc2d4fa74, 32'hc20e8730} /* (4, 8, 7) {real, imag} */,
  {32'h420d9c72, 32'hc2797924} /* (4, 8, 6) {real, imag} */,
  {32'h42e5fea1, 32'h42ebd2ff} /* (4, 8, 5) {real, imag} */,
  {32'h409028c0, 32'hc10a057e} /* (4, 8, 4) {real, imag} */,
  {32'h43181eb1, 32'h4294ea3a} /* (4, 8, 3) {real, imag} */,
  {32'h440843b4, 32'hc2bafe97} /* (4, 8, 2) {real, imag} */,
  {32'hc44c0b48, 32'h42ddaa3a} /* (4, 8, 1) {real, imag} */,
  {32'hc208d678, 32'h00000000} /* (4, 8, 0) {real, imag} */,
  {32'hc455fa23, 32'h42a3454c} /* (4, 7, 31) {real, imag} */,
  {32'h44206f50, 32'h42068963} /* (4, 7, 30) {real, imag} */,
  {32'h437f0584, 32'hc3008de4} /* (4, 7, 29) {real, imag} */,
  {32'h4284f14d, 32'hc24a2d1e} /* (4, 7, 28) {real, imag} */,
  {32'h400513a0, 32'h417aeb14} /* (4, 7, 27) {real, imag} */,
  {32'hc16bab6c, 32'h42bdf560} /* (4, 7, 26) {real, imag} */,
  {32'hc20e89ef, 32'h42730b28} /* (4, 7, 25) {real, imag} */,
  {32'h4113aaa8, 32'hc22fef51} /* (4, 7, 24) {real, imag} */,
  {32'h421079ac, 32'h40a9fb28} /* (4, 7, 23) {real, imag} */,
  {32'hc26ab5ea, 32'hc21d4120} /* (4, 7, 22) {real, imag} */,
  {32'h42b69396, 32'hc239c4ce} /* (4, 7, 21) {real, imag} */,
  {32'hc258682e, 32'h429bf482} /* (4, 7, 20) {real, imag} */,
  {32'hc0037d00, 32'hc14873a8} /* (4, 7, 19) {real, imag} */,
  {32'h42695f75, 32'h3ea6b900} /* (4, 7, 18) {real, imag} */,
  {32'hc19dd4e4, 32'h41cf9870} /* (4, 7, 17) {real, imag} */,
  {32'hc328ab3f, 32'h00000000} /* (4, 7, 16) {real, imag} */,
  {32'hc19dd4e4, 32'hc1cf9870} /* (4, 7, 15) {real, imag} */,
  {32'h42695f75, 32'hbea6b900} /* (4, 7, 14) {real, imag} */,
  {32'hc0037d00, 32'h414873a8} /* (4, 7, 13) {real, imag} */,
  {32'hc258682e, 32'hc29bf482} /* (4, 7, 12) {real, imag} */,
  {32'h42b69396, 32'h4239c4ce} /* (4, 7, 11) {real, imag} */,
  {32'hc26ab5ea, 32'h421d4120} /* (4, 7, 10) {real, imag} */,
  {32'h421079ac, 32'hc0a9fb28} /* (4, 7, 9) {real, imag} */,
  {32'h4113aaa8, 32'h422fef51} /* (4, 7, 8) {real, imag} */,
  {32'hc20e89ef, 32'hc2730b28} /* (4, 7, 7) {real, imag} */,
  {32'hc16bab6c, 32'hc2bdf560} /* (4, 7, 6) {real, imag} */,
  {32'h400513a0, 32'hc17aeb14} /* (4, 7, 5) {real, imag} */,
  {32'h4284f14d, 32'h424a2d1e} /* (4, 7, 4) {real, imag} */,
  {32'h437f0584, 32'h43008de4} /* (4, 7, 3) {real, imag} */,
  {32'h44206f50, 32'hc2068963} /* (4, 7, 2) {real, imag} */,
  {32'hc455fa23, 32'hc2a3454c} /* (4, 7, 1) {real, imag} */,
  {32'h4391810f, 32'h00000000} /* (4, 7, 0) {real, imag} */,
  {32'hc42b9e87, 32'h42f07c51} /* (4, 6, 31) {real, imag} */,
  {32'h43d93cbe, 32'h40b870d0} /* (4, 6, 30) {real, imag} */,
  {32'h433a60f7, 32'h42604f80} /* (4, 6, 29) {real, imag} */,
  {32'h42956467, 32'hc230639d} /* (4, 6, 28) {real, imag} */,
  {32'h418d4508, 32'hc27e6443} /* (4, 6, 27) {real, imag} */,
  {32'h42811cbe, 32'h424023c8} /* (4, 6, 26) {real, imag} */,
  {32'h42cfff9a, 32'hc301abf3} /* (4, 6, 25) {real, imag} */,
  {32'hc229b4db, 32'hc1dd882b} /* (4, 6, 24) {real, imag} */,
  {32'hc29c6cb2, 32'hc2167c36} /* (4, 6, 23) {real, imag} */,
  {32'hc2a7edb0, 32'h424fba97} /* (4, 6, 22) {real, imag} */,
  {32'hc2aff515, 32'hc13a42d0} /* (4, 6, 21) {real, imag} */,
  {32'hc1f6356e, 32'h41e72d79} /* (4, 6, 20) {real, imag} */,
  {32'h428bfd1e, 32'h426a07ef} /* (4, 6, 19) {real, imag} */,
  {32'h4293e0f4, 32'h42b2bf3a} /* (4, 6, 18) {real, imag} */,
  {32'h41bca5d0, 32'h419d114f} /* (4, 6, 17) {real, imag} */,
  {32'hc1de661f, 32'h00000000} /* (4, 6, 16) {real, imag} */,
  {32'h41bca5d0, 32'hc19d114f} /* (4, 6, 15) {real, imag} */,
  {32'h4293e0f4, 32'hc2b2bf3a} /* (4, 6, 14) {real, imag} */,
  {32'h428bfd1e, 32'hc26a07ef} /* (4, 6, 13) {real, imag} */,
  {32'hc1f6356e, 32'hc1e72d79} /* (4, 6, 12) {real, imag} */,
  {32'hc2aff515, 32'h413a42d0} /* (4, 6, 11) {real, imag} */,
  {32'hc2a7edb0, 32'hc24fba97} /* (4, 6, 10) {real, imag} */,
  {32'hc29c6cb2, 32'h42167c36} /* (4, 6, 9) {real, imag} */,
  {32'hc229b4db, 32'h41dd882b} /* (4, 6, 8) {real, imag} */,
  {32'h42cfff9a, 32'h4301abf3} /* (4, 6, 7) {real, imag} */,
  {32'h42811cbe, 32'hc24023c8} /* (4, 6, 6) {real, imag} */,
  {32'h418d4508, 32'h427e6443} /* (4, 6, 5) {real, imag} */,
  {32'h42956467, 32'h4230639d} /* (4, 6, 4) {real, imag} */,
  {32'h433a60f7, 32'hc2604f80} /* (4, 6, 3) {real, imag} */,
  {32'h43d93cbe, 32'hc0b870d0} /* (4, 6, 2) {real, imag} */,
  {32'hc42b9e87, 32'hc2f07c51} /* (4, 6, 1) {real, imag} */,
  {32'h4395be7e, 32'h00000000} /* (4, 6, 0) {real, imag} */,
  {32'hc3a0ee50, 32'h4430aa7a} /* (4, 5, 31) {real, imag} */,
  {32'h430cc474, 32'hc157c73c} /* (4, 5, 30) {real, imag} */,
  {32'h4377bf44, 32'hc27cbe94} /* (4, 5, 29) {real, imag} */,
  {32'h41b9ae80, 32'hc37abb40} /* (4, 5, 28) {real, imag} */,
  {32'h42d43f90, 32'hc1994714} /* (4, 5, 27) {real, imag} */,
  {32'hc219b006, 32'h430197cf} /* (4, 5, 26) {real, imag} */,
  {32'h422aa86c, 32'hc23b3646} /* (4, 5, 25) {real, imag} */,
  {32'hc2081ebc, 32'hc2bbc6c3} /* (4, 5, 24) {real, imag} */,
  {32'h41aa0a36, 32'hc1a8785c} /* (4, 5, 23) {real, imag} */,
  {32'hc1d49294, 32'hc2ca2b98} /* (4, 5, 22) {real, imag} */,
  {32'hc22ba03d, 32'h422db562} /* (4, 5, 21) {real, imag} */,
  {32'hc2aed27a, 32'h404842c0} /* (4, 5, 20) {real, imag} */,
  {32'hc1d603de, 32'hc239a88a} /* (4, 5, 19) {real, imag} */,
  {32'h42b5fb9e, 32'h42574b2b} /* (4, 5, 18) {real, imag} */,
  {32'hc0dd7b89, 32'h422d7dfc} /* (4, 5, 17) {real, imag} */,
  {32'h42c39893, 32'h00000000} /* (4, 5, 16) {real, imag} */,
  {32'hc0dd7b89, 32'hc22d7dfc} /* (4, 5, 15) {real, imag} */,
  {32'h42b5fb9e, 32'hc2574b2b} /* (4, 5, 14) {real, imag} */,
  {32'hc1d603de, 32'h4239a88a} /* (4, 5, 13) {real, imag} */,
  {32'hc2aed27a, 32'hc04842c0} /* (4, 5, 12) {real, imag} */,
  {32'hc22ba03d, 32'hc22db562} /* (4, 5, 11) {real, imag} */,
  {32'hc1d49294, 32'h42ca2b98} /* (4, 5, 10) {real, imag} */,
  {32'h41aa0a36, 32'h41a8785c} /* (4, 5, 9) {real, imag} */,
  {32'hc2081ebc, 32'h42bbc6c3} /* (4, 5, 8) {real, imag} */,
  {32'h422aa86c, 32'h423b3646} /* (4, 5, 7) {real, imag} */,
  {32'hc219b006, 32'hc30197cf} /* (4, 5, 6) {real, imag} */,
  {32'h42d43f90, 32'h41994714} /* (4, 5, 5) {real, imag} */,
  {32'h41b9ae80, 32'h437abb40} /* (4, 5, 4) {real, imag} */,
  {32'h4377bf44, 32'h427cbe94} /* (4, 5, 3) {real, imag} */,
  {32'h430cc474, 32'h4157c73c} /* (4, 5, 2) {real, imag} */,
  {32'hc3a0ee50, 32'hc430aa7a} /* (4, 5, 1) {real, imag} */,
  {32'h4341d8dd, 32'h00000000} /* (4, 5, 0) {real, imag} */,
  {32'hc37cbde3, 32'h445903e8} /* (4, 4, 31) {real, imag} */,
  {32'hc3026e7f, 32'hc34f05e7} /* (4, 4, 30) {real, imag} */,
  {32'h432fedab, 32'hc22583e8} /* (4, 4, 29) {real, imag} */,
  {32'h427d4370, 32'hc38b6a0b} /* (4, 4, 28) {real, imag} */,
  {32'h438bfed5, 32'h423d09bb} /* (4, 4, 27) {real, imag} */,
  {32'h42b0f4fa, 32'hc28f3344} /* (4, 4, 26) {real, imag} */,
  {32'hc1f168d6, 32'hc2f403d3} /* (4, 4, 25) {real, imag} */,
  {32'hc3452a7e, 32'hc1eae17c} /* (4, 4, 24) {real, imag} */,
  {32'hc2359465, 32'h425c68b0} /* (4, 4, 23) {real, imag} */,
  {32'hc1aa6a23, 32'hc214dc7e} /* (4, 4, 22) {real, imag} */,
  {32'h40ea9568, 32'hc2a1ca23} /* (4, 4, 21) {real, imag} */,
  {32'h420538c0, 32'h4221951c} /* (4, 4, 20) {real, imag} */,
  {32'h4264a8ea, 32'h424e3f94} /* (4, 4, 19) {real, imag} */,
  {32'hc29536eb, 32'hc29e2977} /* (4, 4, 18) {real, imag} */,
  {32'hc08d76c4, 32'h410ec06a} /* (4, 4, 17) {real, imag} */,
  {32'hc10b4f5e, 32'h00000000} /* (4, 4, 16) {real, imag} */,
  {32'hc08d76c4, 32'hc10ec06a} /* (4, 4, 15) {real, imag} */,
  {32'hc29536eb, 32'h429e2977} /* (4, 4, 14) {real, imag} */,
  {32'h4264a8ea, 32'hc24e3f94} /* (4, 4, 13) {real, imag} */,
  {32'h420538c0, 32'hc221951c} /* (4, 4, 12) {real, imag} */,
  {32'h40ea9568, 32'h42a1ca23} /* (4, 4, 11) {real, imag} */,
  {32'hc1aa6a23, 32'h4214dc7e} /* (4, 4, 10) {real, imag} */,
  {32'hc2359465, 32'hc25c68b0} /* (4, 4, 9) {real, imag} */,
  {32'hc3452a7e, 32'h41eae17c} /* (4, 4, 8) {real, imag} */,
  {32'hc1f168d6, 32'h42f403d3} /* (4, 4, 7) {real, imag} */,
  {32'h42b0f4fa, 32'h428f3344} /* (4, 4, 6) {real, imag} */,
  {32'h438bfed5, 32'hc23d09bb} /* (4, 4, 5) {real, imag} */,
  {32'h427d4370, 32'h438b6a0b} /* (4, 4, 4) {real, imag} */,
  {32'h432fedab, 32'h422583e8} /* (4, 4, 3) {real, imag} */,
  {32'hc3026e7f, 32'h434f05e7} /* (4, 4, 2) {real, imag} */,
  {32'hc37cbde3, 32'hc45903e8} /* (4, 4, 1) {real, imag} */,
  {32'h435bbf7b, 32'h00000000} /* (4, 4, 0) {real, imag} */,
  {32'hc2d33e40, 32'h4449c635} /* (4, 3, 31) {real, imag} */,
  {32'hc3b0a2ee, 32'hc3a09109} /* (4, 3, 30) {real, imag} */,
  {32'h42e7886a, 32'h429d8ba1} /* (4, 3, 29) {real, imag} */,
  {32'h4251a26e, 32'hc39c01ae} /* (4, 3, 28) {real, imag} */,
  {32'h439f1eea, 32'h42a19293} /* (4, 3, 27) {real, imag} */,
  {32'h430e2cd4, 32'hc30a3358} /* (4, 3, 26) {real, imag} */,
  {32'h42a4bb50, 32'h4235faa8} /* (4, 3, 25) {real, imag} */,
  {32'hc302b846, 32'h426309f5} /* (4, 3, 24) {real, imag} */,
  {32'hc221af9a, 32'hc253b53e} /* (4, 3, 23) {real, imag} */,
  {32'hc17057bf, 32'h42a73662} /* (4, 3, 22) {real, imag} */,
  {32'h4118db7e, 32'hc0197d00} /* (4, 3, 21) {real, imag} */,
  {32'h42258621, 32'hc223314d} /* (4, 3, 20) {real, imag} */,
  {32'h41bf94f8, 32'h40a1a298} /* (4, 3, 19) {real, imag} */,
  {32'h415b2c64, 32'hc2058a46} /* (4, 3, 18) {real, imag} */,
  {32'h421d7f33, 32'hc222af3e} /* (4, 3, 17) {real, imag} */,
  {32'hc14f0c4a, 32'h00000000} /* (4, 3, 16) {real, imag} */,
  {32'h421d7f33, 32'h4222af3e} /* (4, 3, 15) {real, imag} */,
  {32'h415b2c64, 32'h42058a46} /* (4, 3, 14) {real, imag} */,
  {32'h41bf94f8, 32'hc0a1a298} /* (4, 3, 13) {real, imag} */,
  {32'h42258621, 32'h4223314d} /* (4, 3, 12) {real, imag} */,
  {32'h4118db7e, 32'h40197d00} /* (4, 3, 11) {real, imag} */,
  {32'hc17057bf, 32'hc2a73662} /* (4, 3, 10) {real, imag} */,
  {32'hc221af9a, 32'h4253b53e} /* (4, 3, 9) {real, imag} */,
  {32'hc302b846, 32'hc26309f5} /* (4, 3, 8) {real, imag} */,
  {32'h42a4bb50, 32'hc235faa8} /* (4, 3, 7) {real, imag} */,
  {32'h430e2cd4, 32'h430a3358} /* (4, 3, 6) {real, imag} */,
  {32'h439f1eea, 32'hc2a19293} /* (4, 3, 5) {real, imag} */,
  {32'h4251a26e, 32'h439c01ae} /* (4, 3, 4) {real, imag} */,
  {32'h42e7886a, 32'hc29d8ba1} /* (4, 3, 3) {real, imag} */,
  {32'hc3b0a2ee, 32'h43a09109} /* (4, 3, 2) {real, imag} */,
  {32'hc2d33e40, 32'hc449c635} /* (4, 3, 1) {real, imag} */,
  {32'h43e68661, 32'h00000000} /* (4, 3, 0) {real, imag} */,
  {32'hc2c54276, 32'h443d54ac} /* (4, 2, 31) {real, imag} */,
  {32'hc3aebfe1, 32'hc3c56f14} /* (4, 2, 30) {real, imag} */,
  {32'h42dd65d3, 32'h4294792e} /* (4, 2, 29) {real, imag} */,
  {32'h4346066a, 32'hc3ac8e89} /* (4, 2, 28) {real, imag} */,
  {32'h42ad787a, 32'hc259e396} /* (4, 2, 27) {real, imag} */,
  {32'h4203f3fa, 32'h4284bf2d} /* (4, 2, 26) {real, imag} */,
  {32'hc0796950, 32'h424ac0f7} /* (4, 2, 25) {real, imag} */,
  {32'h41f51c06, 32'hc12abd24} /* (4, 2, 24) {real, imag} */,
  {32'h414796ec, 32'h42a2fdbb} /* (4, 2, 23) {real, imag} */,
  {32'hc28f49d6, 32'hc30f8986} /* (4, 2, 22) {real, imag} */,
  {32'h426ff39c, 32'h425dc4ae} /* (4, 2, 21) {real, imag} */,
  {32'hc11cac04, 32'hc1900992} /* (4, 2, 20) {real, imag} */,
  {32'h4306c5b4, 32'hc2a6a6b3} /* (4, 2, 19) {real, imag} */,
  {32'hc219ddf1, 32'hc06f42d0} /* (4, 2, 18) {real, imag} */,
  {32'hc1880eea, 32'hc28639f0} /* (4, 2, 17) {real, imag} */,
  {32'h41bec5c0, 32'h00000000} /* (4, 2, 16) {real, imag} */,
  {32'hc1880eea, 32'h428639f0} /* (4, 2, 15) {real, imag} */,
  {32'hc219ddf1, 32'h406f42d0} /* (4, 2, 14) {real, imag} */,
  {32'h4306c5b4, 32'h42a6a6b3} /* (4, 2, 13) {real, imag} */,
  {32'hc11cac04, 32'h41900992} /* (4, 2, 12) {real, imag} */,
  {32'h426ff39c, 32'hc25dc4ae} /* (4, 2, 11) {real, imag} */,
  {32'hc28f49d6, 32'h430f8986} /* (4, 2, 10) {real, imag} */,
  {32'h414796ec, 32'hc2a2fdbb} /* (4, 2, 9) {real, imag} */,
  {32'h41f51c06, 32'h412abd24} /* (4, 2, 8) {real, imag} */,
  {32'hc0796950, 32'hc24ac0f7} /* (4, 2, 7) {real, imag} */,
  {32'h4203f3fa, 32'hc284bf2d} /* (4, 2, 6) {real, imag} */,
  {32'h42ad787a, 32'h4259e396} /* (4, 2, 5) {real, imag} */,
  {32'h4346066a, 32'h43ac8e89} /* (4, 2, 4) {real, imag} */,
  {32'h42dd65d3, 32'hc294792e} /* (4, 2, 3) {real, imag} */,
  {32'hc3aebfe1, 32'h43c56f14} /* (4, 2, 2) {real, imag} */,
  {32'hc2c54276, 32'hc43d54ac} /* (4, 2, 1) {real, imag} */,
  {32'h44176c58, 32'h00000000} /* (4, 2, 0) {real, imag} */,
  {32'hc23221c0, 32'h442a75e5} /* (4, 1, 31) {real, imag} */,
  {32'hc3483878, 32'hc3e12f36} /* (4, 1, 30) {real, imag} */,
  {32'h4306deac, 32'hc1ab8082} /* (4, 1, 29) {real, imag} */,
  {32'h435236bf, 32'hc34951ce} /* (4, 1, 28) {real, imag} */,
  {32'h435d437c, 32'h4307b2c0} /* (4, 1, 27) {real, imag} */,
  {32'hc1c2d56e, 32'h4143c248} /* (4, 1, 26) {real, imag} */,
  {32'hc1a0201a, 32'h4255830a} /* (4, 1, 25) {real, imag} */,
  {32'hc30c8314, 32'h417f8b0c} /* (4, 1, 24) {real, imag} */,
  {32'hc26a2d9d, 32'hc303f6df} /* (4, 1, 23) {real, imag} */,
  {32'h42dba704, 32'hc2934bb4} /* (4, 1, 22) {real, imag} */,
  {32'hc20aabc5, 32'h418937c4} /* (4, 1, 21) {real, imag} */,
  {32'hc1ac2866, 32'h41c9bf20} /* (4, 1, 20) {real, imag} */,
  {32'h4000a584, 32'hc1f0dfd5} /* (4, 1, 19) {real, imag} */,
  {32'hc24aef48, 32'hc0e7b374} /* (4, 1, 18) {real, imag} */,
  {32'h423061c2, 32'h4260fdec} /* (4, 1, 17) {real, imag} */,
  {32'h422221d8, 32'h00000000} /* (4, 1, 16) {real, imag} */,
  {32'h423061c2, 32'hc260fdec} /* (4, 1, 15) {real, imag} */,
  {32'hc24aef48, 32'h40e7b374} /* (4, 1, 14) {real, imag} */,
  {32'h4000a584, 32'h41f0dfd5} /* (4, 1, 13) {real, imag} */,
  {32'hc1ac2866, 32'hc1c9bf20} /* (4, 1, 12) {real, imag} */,
  {32'hc20aabc5, 32'hc18937c4} /* (4, 1, 11) {real, imag} */,
  {32'h42dba704, 32'h42934bb4} /* (4, 1, 10) {real, imag} */,
  {32'hc26a2d9d, 32'h4303f6df} /* (4, 1, 9) {real, imag} */,
  {32'hc30c8314, 32'hc17f8b0c} /* (4, 1, 8) {real, imag} */,
  {32'hc1a0201a, 32'hc255830a} /* (4, 1, 7) {real, imag} */,
  {32'hc1c2d56e, 32'hc143c248} /* (4, 1, 6) {real, imag} */,
  {32'h435d437c, 32'hc307b2c0} /* (4, 1, 5) {real, imag} */,
  {32'h435236bf, 32'h434951ce} /* (4, 1, 4) {real, imag} */,
  {32'h4306deac, 32'h41ab8082} /* (4, 1, 3) {real, imag} */,
  {32'hc3483878, 32'h43e12f36} /* (4, 1, 2) {real, imag} */,
  {32'hc23221c0, 32'hc42a75e5} /* (4, 1, 1) {real, imag} */,
  {32'h44444fac, 32'h00000000} /* (4, 1, 0) {real, imag} */,
  {32'hc27bf8b8, 32'h43ba1aa6} /* (4, 0, 31) {real, imag} */,
  {32'h419bc570, 32'hc3a8660a} /* (4, 0, 30) {real, imag} */,
  {32'h424a2e52, 32'hc222c478} /* (4, 0, 29) {real, imag} */,
  {32'h428129c8, 32'hc31bb62e} /* (4, 0, 28) {real, imag} */,
  {32'h4355c92e, 32'h42a5c08d} /* (4, 0, 27) {real, imag} */,
  {32'hc05acb08, 32'h3e624680} /* (4, 0, 26) {real, imag} */,
  {32'hc229663b, 32'hc16b1e80} /* (4, 0, 25) {real, imag} */,
  {32'hc2cd60dc, 32'hc18ffd64} /* (4, 0, 24) {real, imag} */,
  {32'hc22d4d1b, 32'hc3057d21} /* (4, 0, 23) {real, imag} */,
  {32'hc0d0494c, 32'hc253f12f} /* (4, 0, 22) {real, imag} */,
  {32'hc26fe052, 32'h42aa142c} /* (4, 0, 21) {real, imag} */,
  {32'h4206ac6a, 32'h41bbbe14} /* (4, 0, 20) {real, imag} */,
  {32'hc224dffc, 32'h40516cc4} /* (4, 0, 19) {real, imag} */,
  {32'h3fb9c900, 32'hc202ed28} /* (4, 0, 18) {real, imag} */,
  {32'h418ede9a, 32'h421df923} /* (4, 0, 17) {real, imag} */,
  {32'h41c5448c, 32'h00000000} /* (4, 0, 16) {real, imag} */,
  {32'h418ede9a, 32'hc21df923} /* (4, 0, 15) {real, imag} */,
  {32'h3fb9c900, 32'h4202ed28} /* (4, 0, 14) {real, imag} */,
  {32'hc224dffc, 32'hc0516cc4} /* (4, 0, 13) {real, imag} */,
  {32'h4206ac6a, 32'hc1bbbe14} /* (4, 0, 12) {real, imag} */,
  {32'hc26fe052, 32'hc2aa142c} /* (4, 0, 11) {real, imag} */,
  {32'hc0d0494c, 32'h4253f12f} /* (4, 0, 10) {real, imag} */,
  {32'hc22d4d1b, 32'h43057d21} /* (4, 0, 9) {real, imag} */,
  {32'hc2cd60dc, 32'h418ffd64} /* (4, 0, 8) {real, imag} */,
  {32'hc229663b, 32'h416b1e80} /* (4, 0, 7) {real, imag} */,
  {32'hc05acb08, 32'hbe624680} /* (4, 0, 6) {real, imag} */,
  {32'h4355c92e, 32'hc2a5c08d} /* (4, 0, 5) {real, imag} */,
  {32'h428129c8, 32'h431bb62e} /* (4, 0, 4) {real, imag} */,
  {32'h424a2e52, 32'h4222c478} /* (4, 0, 3) {real, imag} */,
  {32'h419bc570, 32'h43a8660a} /* (4, 0, 2) {real, imag} */,
  {32'hc27bf8b8, 32'hc3ba1aa6} /* (4, 0, 1) {real, imag} */,
  {32'h4467531c, 32'h00000000} /* (4, 0, 0) {real, imag} */,
  {32'hc464e8e5, 32'h43d8b39f} /* (3, 31, 31) {real, imag} */,
  {32'h43eaa161, 32'hc38238fd} /* (3, 31, 30) {real, imag} */,
  {32'h42d16516, 32'hc18f752c} /* (3, 31, 29) {real, imag} */,
  {32'hc30246a0, 32'hc30d597e} /* (3, 31, 28) {real, imag} */,
  {32'h432dcc56, 32'hc2d3e0e9} /* (3, 31, 27) {real, imag} */,
  {32'hc1b2a054, 32'hc2a723ae} /* (3, 31, 26) {real, imag} */,
  {32'h40a64d80, 32'h412a9c0c} /* (3, 31, 25) {real, imag} */,
  {32'hc277a12a, 32'hc209419c} /* (3, 31, 24) {real, imag} */,
  {32'h427a42f8, 32'hc1b30842} /* (3, 31, 23) {real, imag} */,
  {32'hc00365a0, 32'h42638480} /* (3, 31, 22) {real, imag} */,
  {32'hc1e3daff, 32'hc2190182} /* (3, 31, 21) {real, imag} */,
  {32'h41a1346f, 32'h41d5e72d} /* (3, 31, 20) {real, imag} */,
  {32'hc2adc98e, 32'hc27d84f2} /* (3, 31, 19) {real, imag} */,
  {32'h41b91514, 32'h420c226b} /* (3, 31, 18) {real, imag} */,
  {32'h40f26278, 32'h41ea1c53} /* (3, 31, 17) {real, imag} */,
  {32'h40926c48, 32'h00000000} /* (3, 31, 16) {real, imag} */,
  {32'h40f26278, 32'hc1ea1c53} /* (3, 31, 15) {real, imag} */,
  {32'h41b91514, 32'hc20c226b} /* (3, 31, 14) {real, imag} */,
  {32'hc2adc98e, 32'h427d84f2} /* (3, 31, 13) {real, imag} */,
  {32'h41a1346f, 32'hc1d5e72d} /* (3, 31, 12) {real, imag} */,
  {32'hc1e3daff, 32'h42190182} /* (3, 31, 11) {real, imag} */,
  {32'hc00365a0, 32'hc2638480} /* (3, 31, 10) {real, imag} */,
  {32'h427a42f8, 32'h41b30842} /* (3, 31, 9) {real, imag} */,
  {32'hc277a12a, 32'h4209419c} /* (3, 31, 8) {real, imag} */,
  {32'h40a64d80, 32'hc12a9c0c} /* (3, 31, 7) {real, imag} */,
  {32'hc1b2a054, 32'h42a723ae} /* (3, 31, 6) {real, imag} */,
  {32'h432dcc56, 32'h42d3e0e9} /* (3, 31, 5) {real, imag} */,
  {32'hc30246a0, 32'h430d597e} /* (3, 31, 4) {real, imag} */,
  {32'h42d16516, 32'h418f752c} /* (3, 31, 3) {real, imag} */,
  {32'h43eaa161, 32'h438238fd} /* (3, 31, 2) {real, imag} */,
  {32'hc464e8e5, 32'hc3d8b39f} /* (3, 31, 1) {real, imag} */,
  {32'h41d7d49e, 32'h00000000} /* (3, 31, 0) {real, imag} */,
  {32'hc4983df4, 32'h4386d55a} /* (3, 30, 31) {real, imag} */,
  {32'h4457da4c, 32'hc353431e} /* (3, 30, 30) {real, imag} */,
  {32'h43463afb, 32'hc1b69f1c} /* (3, 30, 29) {real, imag} */,
  {32'hc31baa64, 32'hc2848804} /* (3, 30, 28) {real, imag} */,
  {32'h437563da, 32'hc359921c} /* (3, 30, 27) {real, imag} */,
  {32'h40e25a40, 32'h4109adc0} /* (3, 30, 26) {real, imag} */,
  {32'hc19cbeb6, 32'h428632f2} /* (3, 30, 25) {real, imag} */,
  {32'h42c11a11, 32'hc18f0f85} /* (3, 30, 24) {real, imag} */,
  {32'h425f6dc4, 32'h4317cb78} /* (3, 30, 23) {real, imag} */,
  {32'hc070a2a8, 32'h402d6140} /* (3, 30, 22) {real, imag} */,
  {32'hc1cd7c04, 32'hc29b9352} /* (3, 30, 21) {real, imag} */,
  {32'h42778514, 32'h417b58f6} /* (3, 30, 20) {real, imag} */,
  {32'h428c57e9, 32'h4251aafc} /* (3, 30, 19) {real, imag} */,
  {32'h41e8059c, 32'h41521cfc} /* (3, 30, 18) {real, imag} */,
  {32'hc09f8030, 32'h42212b86} /* (3, 30, 17) {real, imag} */,
  {32'hc1f60225, 32'h00000000} /* (3, 30, 16) {real, imag} */,
  {32'hc09f8030, 32'hc2212b86} /* (3, 30, 15) {real, imag} */,
  {32'h41e8059c, 32'hc1521cfc} /* (3, 30, 14) {real, imag} */,
  {32'h428c57e9, 32'hc251aafc} /* (3, 30, 13) {real, imag} */,
  {32'h42778514, 32'hc17b58f6} /* (3, 30, 12) {real, imag} */,
  {32'hc1cd7c04, 32'h429b9352} /* (3, 30, 11) {real, imag} */,
  {32'hc070a2a8, 32'hc02d6140} /* (3, 30, 10) {real, imag} */,
  {32'h425f6dc4, 32'hc317cb78} /* (3, 30, 9) {real, imag} */,
  {32'h42c11a11, 32'h418f0f85} /* (3, 30, 8) {real, imag} */,
  {32'hc19cbeb6, 32'hc28632f2} /* (3, 30, 7) {real, imag} */,
  {32'h40e25a40, 32'hc109adc0} /* (3, 30, 6) {real, imag} */,
  {32'h437563da, 32'h4359921c} /* (3, 30, 5) {real, imag} */,
  {32'hc31baa64, 32'h42848804} /* (3, 30, 4) {real, imag} */,
  {32'h43463afb, 32'h41b69f1c} /* (3, 30, 3) {real, imag} */,
  {32'h4457da4c, 32'h4353431e} /* (3, 30, 2) {real, imag} */,
  {32'hc4983df4, 32'hc386d55a} /* (3, 30, 1) {real, imag} */,
  {32'hc30eb332, 32'h00000000} /* (3, 30, 0) {real, imag} */,
  {32'hc4bd00cc, 32'h435842d4} /* (3, 29, 31) {real, imag} */,
  {32'h4472b250, 32'hc23b4328} /* (3, 29, 30) {real, imag} */,
  {32'h4362d306, 32'hc30d97c6} /* (3, 29, 29) {real, imag} */,
  {32'hc35d244b, 32'h42ffad80} /* (3, 29, 28) {real, imag} */,
  {32'h438449e0, 32'hc32054c2} /* (3, 29, 27) {real, imag} */,
  {32'h429b8a0d, 32'h4333170f} /* (3, 29, 26) {real, imag} */,
  {32'hc2bdf93e, 32'h42d9092a} /* (3, 29, 25) {real, imag} */,
  {32'h42db7598, 32'hc2b5def2} /* (3, 29, 24) {real, imag} */,
  {32'hc2ac9462, 32'h4328aa4d} /* (3, 29, 23) {real, imag} */,
  {32'hc17a43e6, 32'hc2972daf} /* (3, 29, 22) {real, imag} */,
  {32'h42df393c, 32'hc2e00074} /* (3, 29, 21) {real, imag} */,
  {32'h41fa2d05, 32'hc1b4b24b} /* (3, 29, 20) {real, imag} */,
  {32'h41baf6b6, 32'hc2aa9ae8} /* (3, 29, 19) {real, imag} */,
  {32'hc20af8d4, 32'h42939178} /* (3, 29, 18) {real, imag} */,
  {32'h42085812, 32'hc13a4b5c} /* (3, 29, 17) {real, imag} */,
  {32'h423092ee, 32'h00000000} /* (3, 29, 16) {real, imag} */,
  {32'h42085812, 32'h413a4b5c} /* (3, 29, 15) {real, imag} */,
  {32'hc20af8d4, 32'hc2939178} /* (3, 29, 14) {real, imag} */,
  {32'h41baf6b6, 32'h42aa9ae8} /* (3, 29, 13) {real, imag} */,
  {32'h41fa2d05, 32'h41b4b24b} /* (3, 29, 12) {real, imag} */,
  {32'h42df393c, 32'h42e00074} /* (3, 29, 11) {real, imag} */,
  {32'hc17a43e6, 32'h42972daf} /* (3, 29, 10) {real, imag} */,
  {32'hc2ac9462, 32'hc328aa4d} /* (3, 29, 9) {real, imag} */,
  {32'h42db7598, 32'h42b5def2} /* (3, 29, 8) {real, imag} */,
  {32'hc2bdf93e, 32'hc2d9092a} /* (3, 29, 7) {real, imag} */,
  {32'h429b8a0d, 32'hc333170f} /* (3, 29, 6) {real, imag} */,
  {32'h438449e0, 32'h432054c2} /* (3, 29, 5) {real, imag} */,
  {32'hc35d244b, 32'hc2ffad80} /* (3, 29, 4) {real, imag} */,
  {32'h4362d306, 32'h430d97c6} /* (3, 29, 3) {real, imag} */,
  {32'h4472b250, 32'h423b4328} /* (3, 29, 2) {real, imag} */,
  {32'hc4bd00cc, 32'hc35842d4} /* (3, 29, 1) {real, imag} */,
  {32'hc25f7230, 32'h00000000} /* (3, 29, 0) {real, imag} */,
  {32'hc4c60a33, 32'h435154b4} /* (3, 28, 31) {real, imag} */,
  {32'h446e40ac, 32'hc24e5490} /* (3, 28, 30) {real, imag} */,
  {32'h4307166b, 32'hc2a4d3f2} /* (3, 28, 29) {real, imag} */,
  {32'hc2c47b8a, 32'h4243be18} /* (3, 28, 28) {real, imag} */,
  {32'h4378983f, 32'hc340c61a} /* (3, 28, 27) {real, imag} */,
  {32'h422ab758, 32'hc21c5139} /* (3, 28, 26) {real, imag} */,
  {32'hc30c9add, 32'h42b233f3} /* (3, 28, 25) {real, imag} */,
  {32'h42a0e498, 32'hc1be1a17} /* (3, 28, 24) {real, imag} */,
  {32'hc2b898f0, 32'h427ed28d} /* (3, 28, 23) {real, imag} */,
  {32'h429eb91b, 32'h41274fbc} /* (3, 28, 22) {real, imag} */,
  {32'h429f8baa, 32'hc2a8f441} /* (3, 28, 21) {real, imag} */,
  {32'hc29852e0, 32'h41561e40} /* (3, 28, 20) {real, imag} */,
  {32'hc2a02b6a, 32'hc27f8bd8} /* (3, 28, 19) {real, imag} */,
  {32'hc1ca87a2, 32'h427e4d03} /* (3, 28, 18) {real, imag} */,
  {32'hc19752c4, 32'hc2580c38} /* (3, 28, 17) {real, imag} */,
  {32'h4299997a, 32'h00000000} /* (3, 28, 16) {real, imag} */,
  {32'hc19752c4, 32'h42580c38} /* (3, 28, 15) {real, imag} */,
  {32'hc1ca87a2, 32'hc27e4d03} /* (3, 28, 14) {real, imag} */,
  {32'hc2a02b6a, 32'h427f8bd8} /* (3, 28, 13) {real, imag} */,
  {32'hc29852e0, 32'hc1561e40} /* (3, 28, 12) {real, imag} */,
  {32'h429f8baa, 32'h42a8f441} /* (3, 28, 11) {real, imag} */,
  {32'h429eb91b, 32'hc1274fbc} /* (3, 28, 10) {real, imag} */,
  {32'hc2b898f0, 32'hc27ed28d} /* (3, 28, 9) {real, imag} */,
  {32'h42a0e498, 32'h41be1a17} /* (3, 28, 8) {real, imag} */,
  {32'hc30c9add, 32'hc2b233f3} /* (3, 28, 7) {real, imag} */,
  {32'h422ab758, 32'h421c5139} /* (3, 28, 6) {real, imag} */,
  {32'h4378983f, 32'h4340c61a} /* (3, 28, 5) {real, imag} */,
  {32'hc2c47b8a, 32'hc243be18} /* (3, 28, 4) {real, imag} */,
  {32'h4307166b, 32'h42a4d3f2} /* (3, 28, 3) {real, imag} */,
  {32'h446e40ac, 32'h424e5490} /* (3, 28, 2) {real, imag} */,
  {32'hc4c60a33, 32'hc35154b4} /* (3, 28, 1) {real, imag} */,
  {32'hc30a229e, 32'h00000000} /* (3, 28, 0) {real, imag} */,
  {32'hc4c9d310, 32'h435365fc} /* (3, 27, 31) {real, imag} */,
  {32'h446699d0, 32'hc30c634a} /* (3, 27, 30) {real, imag} */,
  {32'h42e74080, 32'hc338f329} /* (3, 27, 29) {real, imag} */,
  {32'hc3709a96, 32'h41b0a880} /* (3, 27, 28) {real, imag} */,
  {32'h439e1683, 32'hc2b9de13} /* (3, 27, 27) {real, imag} */,
  {32'hc2a52ffb, 32'h409d7162} /* (3, 27, 26) {real, imag} */,
  {32'hc200996a, 32'hc1529380} /* (3, 27, 25) {real, imag} */,
  {32'h42f3aa50, 32'hc1cb8dba} /* (3, 27, 24) {real, imag} */,
  {32'h40e57340, 32'hc15b1bba} /* (3, 27, 23) {real, imag} */,
  {32'hc25be0ca, 32'hc26601e4} /* (3, 27, 22) {real, imag} */,
  {32'h40748b90, 32'hc1a6d175} /* (3, 27, 21) {real, imag} */,
  {32'h4299027f, 32'h40d178ac} /* (3, 27, 20) {real, imag} */,
  {32'h41c357c6, 32'hc2423ca3} /* (3, 27, 19) {real, imag} */,
  {32'h4247b34c, 32'hc18fec66} /* (3, 27, 18) {real, imag} */,
  {32'h430658ff, 32'h42377bb4} /* (3, 27, 17) {real, imag} */,
  {32'hc24cd1be, 32'h00000000} /* (3, 27, 16) {real, imag} */,
  {32'h430658ff, 32'hc2377bb4} /* (3, 27, 15) {real, imag} */,
  {32'h4247b34c, 32'h418fec66} /* (3, 27, 14) {real, imag} */,
  {32'h41c357c6, 32'h42423ca3} /* (3, 27, 13) {real, imag} */,
  {32'h4299027f, 32'hc0d178ac} /* (3, 27, 12) {real, imag} */,
  {32'h40748b90, 32'h41a6d175} /* (3, 27, 11) {real, imag} */,
  {32'hc25be0ca, 32'h426601e4} /* (3, 27, 10) {real, imag} */,
  {32'h40e57340, 32'h415b1bba} /* (3, 27, 9) {real, imag} */,
  {32'h42f3aa50, 32'h41cb8dba} /* (3, 27, 8) {real, imag} */,
  {32'hc200996a, 32'h41529380} /* (3, 27, 7) {real, imag} */,
  {32'hc2a52ffb, 32'hc09d7162} /* (3, 27, 6) {real, imag} */,
  {32'h439e1683, 32'h42b9de13} /* (3, 27, 5) {real, imag} */,
  {32'hc3709a96, 32'hc1b0a880} /* (3, 27, 4) {real, imag} */,
  {32'h42e74080, 32'h4338f329} /* (3, 27, 3) {real, imag} */,
  {32'h446699d0, 32'h430c634a} /* (3, 27, 2) {real, imag} */,
  {32'hc4c9d310, 32'hc35365fc} /* (3, 27, 1) {real, imag} */,
  {32'hc3642319, 32'h00000000} /* (3, 27, 0) {real, imag} */,
  {32'hc4d83ec4, 32'h435de436} /* (3, 26, 31) {real, imag} */,
  {32'h4478e066, 32'hc266a843} /* (3, 26, 30) {real, imag} */,
  {32'h42bfee93, 32'hc347d18a} /* (3, 26, 29) {real, imag} */,
  {32'hc39c720a, 32'h423e5144} /* (3, 26, 28) {real, imag} */,
  {32'h43492139, 32'hc15ad504} /* (3, 26, 27) {real, imag} */,
  {32'h42617054, 32'hc2c52d30} /* (3, 26, 26) {real, imag} */,
  {32'hc2613278, 32'h41096d74} /* (3, 26, 25) {real, imag} */,
  {32'h4228939b, 32'hc2c6f64a} /* (3, 26, 24) {real, imag} */,
  {32'h42a881f0, 32'hc286f9f6} /* (3, 26, 23) {real, imag} */,
  {32'h41192288, 32'h41487a1c} /* (3, 26, 22) {real, imag} */,
  {32'h42732255, 32'h424a39f3} /* (3, 26, 21) {real, imag} */,
  {32'hc2fcb133, 32'h41fef283} /* (3, 26, 20) {real, imag} */,
  {32'h410e4e88, 32'h4285a1e1} /* (3, 26, 19) {real, imag} */,
  {32'hc25cca30, 32'hbe4c1c80} /* (3, 26, 18) {real, imag} */,
  {32'h4203b766, 32'h418f1328} /* (3, 26, 17) {real, imag} */,
  {32'h41cff680, 32'h00000000} /* (3, 26, 16) {real, imag} */,
  {32'h4203b766, 32'hc18f1328} /* (3, 26, 15) {real, imag} */,
  {32'hc25cca30, 32'h3e4c1c80} /* (3, 26, 14) {real, imag} */,
  {32'h410e4e88, 32'hc285a1e1} /* (3, 26, 13) {real, imag} */,
  {32'hc2fcb133, 32'hc1fef283} /* (3, 26, 12) {real, imag} */,
  {32'h42732255, 32'hc24a39f3} /* (3, 26, 11) {real, imag} */,
  {32'h41192288, 32'hc1487a1c} /* (3, 26, 10) {real, imag} */,
  {32'h42a881f0, 32'h4286f9f6} /* (3, 26, 9) {real, imag} */,
  {32'h4228939b, 32'h42c6f64a} /* (3, 26, 8) {real, imag} */,
  {32'hc2613278, 32'hc1096d74} /* (3, 26, 7) {real, imag} */,
  {32'h42617054, 32'h42c52d30} /* (3, 26, 6) {real, imag} */,
  {32'h43492139, 32'h415ad504} /* (3, 26, 5) {real, imag} */,
  {32'hc39c720a, 32'hc23e5144} /* (3, 26, 4) {real, imag} */,
  {32'h42bfee93, 32'h4347d18a} /* (3, 26, 3) {real, imag} */,
  {32'h4478e066, 32'h4266a843} /* (3, 26, 2) {real, imag} */,
  {32'hc4d83ec4, 32'hc35de436} /* (3, 26, 1) {real, imag} */,
  {32'hc3236832, 32'h00000000} /* (3, 26, 0) {real, imag} */,
  {32'hc4ede8f4, 32'h433fbcd6} /* (3, 25, 31) {real, imag} */,
  {32'h44812c05, 32'h41bb38a0} /* (3, 25, 30) {real, imag} */,
  {32'h42d32e56, 32'hc307a146} /* (3, 25, 29) {real, imag} */,
  {32'hc347106c, 32'h41f149f4} /* (3, 25, 28) {real, imag} */,
  {32'h431e3a0e, 32'hc32c0cad} /* (3, 25, 27) {real, imag} */,
  {32'h3fc1e6a0, 32'hc2c32ee0} /* (3, 25, 26) {real, imag} */,
  {32'hc2e919e4, 32'h424a8a59} /* (3, 25, 25) {real, imag} */,
  {32'h420b5d14, 32'hc2afcd1f} /* (3, 25, 24) {real, imag} */,
  {32'h4295f0de, 32'hc1ca3ede} /* (3, 25, 23) {real, imag} */,
  {32'hc18d4860, 32'hc1bb3a96} /* (3, 25, 22) {real, imag} */,
  {32'h42886f5e, 32'hc12f97d8} /* (3, 25, 21) {real, imag} */,
  {32'hc223cc10, 32'h422221d9} /* (3, 25, 20) {real, imag} */,
  {32'h4281c768, 32'h423881c7} /* (3, 25, 19) {real, imag} */,
  {32'h41165097, 32'h4252cedd} /* (3, 25, 18) {real, imag} */,
  {32'hc21646fc, 32'hc29c29c6} /* (3, 25, 17) {real, imag} */,
  {32'hc11dfd8a, 32'h00000000} /* (3, 25, 16) {real, imag} */,
  {32'hc21646fc, 32'h429c29c6} /* (3, 25, 15) {real, imag} */,
  {32'h41165097, 32'hc252cedd} /* (3, 25, 14) {real, imag} */,
  {32'h4281c768, 32'hc23881c7} /* (3, 25, 13) {real, imag} */,
  {32'hc223cc10, 32'hc22221d9} /* (3, 25, 12) {real, imag} */,
  {32'h42886f5e, 32'h412f97d8} /* (3, 25, 11) {real, imag} */,
  {32'hc18d4860, 32'h41bb3a96} /* (3, 25, 10) {real, imag} */,
  {32'h4295f0de, 32'h41ca3ede} /* (3, 25, 9) {real, imag} */,
  {32'h420b5d14, 32'h42afcd1f} /* (3, 25, 8) {real, imag} */,
  {32'hc2e919e4, 32'hc24a8a59} /* (3, 25, 7) {real, imag} */,
  {32'h3fc1e6a0, 32'h42c32ee0} /* (3, 25, 6) {real, imag} */,
  {32'h431e3a0e, 32'h432c0cad} /* (3, 25, 5) {real, imag} */,
  {32'hc347106c, 32'hc1f149f4} /* (3, 25, 4) {real, imag} */,
  {32'h42d32e56, 32'h4307a146} /* (3, 25, 3) {real, imag} */,
  {32'h44812c05, 32'hc1bb38a0} /* (3, 25, 2) {real, imag} */,
  {32'hc4ede8f4, 32'hc33fbcd6} /* (3, 25, 1) {real, imag} */,
  {32'hc39b0aa2, 32'h00000000} /* (3, 25, 0) {real, imag} */,
  {32'hc4edb06b, 32'h43511e32} /* (3, 24, 31) {real, imag} */,
  {32'h4466a370, 32'h41b6199e} /* (3, 24, 30) {real, imag} */,
  {32'h420b2e12, 32'hc1cb1bfc} /* (3, 24, 29) {real, imag} */,
  {32'hc37cba0e, 32'h412e56cc} /* (3, 24, 28) {real, imag} */,
  {32'h4344bbfb, 32'hc2d0d414} /* (3, 24, 27) {real, imag} */,
  {32'h428be9ac, 32'hc2523243} /* (3, 24, 26) {real, imag} */,
  {32'hc231a31e, 32'hc1651a56} /* (3, 24, 25) {real, imag} */,
  {32'hc0dc4d2c, 32'hc2b60d2c} /* (3, 24, 24) {real, imag} */,
  {32'h4243f84c, 32'h41977534} /* (3, 24, 23) {real, imag} */,
  {32'hc2bbcd6c, 32'h42ae5dc5} /* (3, 24, 22) {real, imag} */,
  {32'h42d7fe55, 32'h41737994} /* (3, 24, 21) {real, imag} */,
  {32'h41736e20, 32'hc1e90599} /* (3, 24, 20) {real, imag} */,
  {32'hc0a1056c, 32'hc35541de} /* (3, 24, 19) {real, imag} */,
  {32'hc221a9ed, 32'hc1536e5a} /* (3, 24, 18) {real, imag} */,
  {32'hc306af85, 32'hc0c66b97} /* (3, 24, 17) {real, imag} */,
  {32'h4045d0ac, 32'h00000000} /* (3, 24, 16) {real, imag} */,
  {32'hc306af85, 32'h40c66b97} /* (3, 24, 15) {real, imag} */,
  {32'hc221a9ed, 32'h41536e5a} /* (3, 24, 14) {real, imag} */,
  {32'hc0a1056c, 32'h435541de} /* (3, 24, 13) {real, imag} */,
  {32'h41736e20, 32'h41e90599} /* (3, 24, 12) {real, imag} */,
  {32'h42d7fe55, 32'hc1737994} /* (3, 24, 11) {real, imag} */,
  {32'hc2bbcd6c, 32'hc2ae5dc5} /* (3, 24, 10) {real, imag} */,
  {32'h4243f84c, 32'hc1977534} /* (3, 24, 9) {real, imag} */,
  {32'hc0dc4d2c, 32'h42b60d2c} /* (3, 24, 8) {real, imag} */,
  {32'hc231a31e, 32'h41651a56} /* (3, 24, 7) {real, imag} */,
  {32'h428be9ac, 32'h42523243} /* (3, 24, 6) {real, imag} */,
  {32'h4344bbfb, 32'h42d0d414} /* (3, 24, 5) {real, imag} */,
  {32'hc37cba0e, 32'hc12e56cc} /* (3, 24, 4) {real, imag} */,
  {32'h420b2e12, 32'h41cb1bfc} /* (3, 24, 3) {real, imag} */,
  {32'h4466a370, 32'hc1b6199e} /* (3, 24, 2) {real, imag} */,
  {32'hc4edb06b, 32'hc3511e32} /* (3, 24, 1) {real, imag} */,
  {32'hc3d3bd76, 32'h00000000} /* (3, 24, 0) {real, imag} */,
  {32'hc4d769aa, 32'h4306e386} /* (3, 23, 31) {real, imag} */,
  {32'h442debbf, 32'hc22ab350} /* (3, 23, 30) {real, imag} */,
  {32'h42d8bca6, 32'h414571d6} /* (3, 23, 29) {real, imag} */,
  {32'hc33b26d9, 32'hc29f1b27} /* (3, 23, 28) {real, imag} */,
  {32'h4379f7a6, 32'hc3202de2} /* (3, 23, 27) {real, imag} */,
  {32'h3fac2760, 32'hc0411760} /* (3, 23, 26) {real, imag} */,
  {32'hc000e140, 32'h4266b118} /* (3, 23, 25) {real, imag} */,
  {32'h42950894, 32'h418b97b2} /* (3, 23, 24) {real, imag} */,
  {32'h412b8ce0, 32'h426792ae} /* (3, 23, 23) {real, imag} */,
  {32'hc234cc56, 32'h42ded8f5} /* (3, 23, 22) {real, imag} */,
  {32'h4223ae14, 32'hc1b461e2} /* (3, 23, 21) {real, imag} */,
  {32'hc291f9d5, 32'hc11e07e4} /* (3, 23, 20) {real, imag} */,
  {32'hc2e87109, 32'hc1923980} /* (3, 23, 19) {real, imag} */,
  {32'h4250d4e0, 32'hc23d2233} /* (3, 23, 18) {real, imag} */,
  {32'h423d9566, 32'hc207efa2} /* (3, 23, 17) {real, imag} */,
  {32'h42046944, 32'h00000000} /* (3, 23, 16) {real, imag} */,
  {32'h423d9566, 32'h4207efa2} /* (3, 23, 15) {real, imag} */,
  {32'h4250d4e0, 32'h423d2233} /* (3, 23, 14) {real, imag} */,
  {32'hc2e87109, 32'h41923980} /* (3, 23, 13) {real, imag} */,
  {32'hc291f9d5, 32'h411e07e4} /* (3, 23, 12) {real, imag} */,
  {32'h4223ae14, 32'h41b461e2} /* (3, 23, 11) {real, imag} */,
  {32'hc234cc56, 32'hc2ded8f5} /* (3, 23, 10) {real, imag} */,
  {32'h412b8ce0, 32'hc26792ae} /* (3, 23, 9) {real, imag} */,
  {32'h42950894, 32'hc18b97b2} /* (3, 23, 8) {real, imag} */,
  {32'hc000e140, 32'hc266b118} /* (3, 23, 7) {real, imag} */,
  {32'h3fac2760, 32'h40411760} /* (3, 23, 6) {real, imag} */,
  {32'h4379f7a6, 32'h43202de2} /* (3, 23, 5) {real, imag} */,
  {32'hc33b26d9, 32'h429f1b27} /* (3, 23, 4) {real, imag} */,
  {32'h42d8bca6, 32'hc14571d6} /* (3, 23, 3) {real, imag} */,
  {32'h442debbf, 32'h422ab350} /* (3, 23, 2) {real, imag} */,
  {32'hc4d769aa, 32'hc306e386} /* (3, 23, 1) {real, imag} */,
  {32'hc3c0857e, 32'h00000000} /* (3, 23, 0) {real, imag} */,
  {32'hc4aa1683, 32'h40cad910} /* (3, 22, 31) {real, imag} */,
  {32'h43f2f46e, 32'h4251b955} /* (3, 22, 30) {real, imag} */,
  {32'h42fd9ae9, 32'h42caa426} /* (3, 22, 29) {real, imag} */,
  {32'hc2b35828, 32'hc28e3f91} /* (3, 22, 28) {real, imag} */,
  {32'h4327262e, 32'hc30455d6} /* (3, 22, 27) {real, imag} */,
  {32'hc1ab80d0, 32'hc14ff440} /* (3, 22, 26) {real, imag} */,
  {32'h425dd04c, 32'hc28a31fc} /* (3, 22, 25) {real, imag} */,
  {32'h423e8e48, 32'h42586b4d} /* (3, 22, 24) {real, imag} */,
  {32'h42e7374e, 32'hc2e43646} /* (3, 22, 23) {real, imag} */,
  {32'h4268c785, 32'hc112499f} /* (3, 22, 22) {real, imag} */,
  {32'hc0d73928, 32'hc299e9e0} /* (3, 22, 21) {real, imag} */,
  {32'h3fc1e1c0, 32'h429a1f6c} /* (3, 22, 20) {real, imag} */,
  {32'hc05f4b60, 32'h429d80d9} /* (3, 22, 19) {real, imag} */,
  {32'hc28edf87, 32'hc21f8c50} /* (3, 22, 18) {real, imag} */,
  {32'h41b077c0, 32'hc2a3c962} /* (3, 22, 17) {real, imag} */,
  {32'h41b3e946, 32'h00000000} /* (3, 22, 16) {real, imag} */,
  {32'h41b077c0, 32'h42a3c962} /* (3, 22, 15) {real, imag} */,
  {32'hc28edf87, 32'h421f8c50} /* (3, 22, 14) {real, imag} */,
  {32'hc05f4b60, 32'hc29d80d9} /* (3, 22, 13) {real, imag} */,
  {32'h3fc1e1c0, 32'hc29a1f6c} /* (3, 22, 12) {real, imag} */,
  {32'hc0d73928, 32'h4299e9e0} /* (3, 22, 11) {real, imag} */,
  {32'h4268c785, 32'h4112499f} /* (3, 22, 10) {real, imag} */,
  {32'h42e7374e, 32'h42e43646} /* (3, 22, 9) {real, imag} */,
  {32'h423e8e48, 32'hc2586b4d} /* (3, 22, 8) {real, imag} */,
  {32'h425dd04c, 32'h428a31fc} /* (3, 22, 7) {real, imag} */,
  {32'hc1ab80d0, 32'h414ff440} /* (3, 22, 6) {real, imag} */,
  {32'h4327262e, 32'h430455d6} /* (3, 22, 5) {real, imag} */,
  {32'hc2b35828, 32'h428e3f91} /* (3, 22, 4) {real, imag} */,
  {32'h42fd9ae9, 32'hc2caa426} /* (3, 22, 3) {real, imag} */,
  {32'h43f2f46e, 32'hc251b955} /* (3, 22, 2) {real, imag} */,
  {32'hc4aa1683, 32'hc0cad910} /* (3, 22, 1) {real, imag} */,
  {32'hc3b6df4d, 32'h00000000} /* (3, 22, 0) {real, imag} */,
  {32'hc3dbf8a2, 32'hc32e74f4} /* (3, 21, 31) {real, imag} */,
  {32'h43202238, 32'hc2064858} /* (3, 21, 30) {real, imag} */,
  {32'hc281a59e, 32'hc247b68f} /* (3, 21, 29) {real, imag} */,
  {32'h4263dc2e, 32'hc2d23f48} /* (3, 21, 28) {real, imag} */,
  {32'h4295ad7c, 32'hc3003f30} /* (3, 21, 27) {real, imag} */,
  {32'hc20e735f, 32'h428790fd} /* (3, 21, 26) {real, imag} */,
  {32'hc2c17232, 32'h428f5583} /* (3, 21, 25) {real, imag} */,
  {32'h3fa72650, 32'h42939d9a} /* (3, 21, 24) {real, imag} */,
  {32'h42cb74d7, 32'hc1b344a4} /* (3, 21, 23) {real, imag} */,
  {32'h426ae4d5, 32'h4215a894} /* (3, 21, 22) {real, imag} */,
  {32'hc2b92c74, 32'hc0071d10} /* (3, 21, 21) {real, imag} */,
  {32'h420ddc2a, 32'hc1c51581} /* (3, 21, 20) {real, imag} */,
  {32'hc199ab76, 32'hc276a5ca} /* (3, 21, 19) {real, imag} */,
  {32'hc12c2db9, 32'hc167f92d} /* (3, 21, 18) {real, imag} */,
  {32'hc1f38768, 32'h41742a9b} /* (3, 21, 17) {real, imag} */,
  {32'h41b813c4, 32'h00000000} /* (3, 21, 16) {real, imag} */,
  {32'hc1f38768, 32'hc1742a9b} /* (3, 21, 15) {real, imag} */,
  {32'hc12c2db9, 32'h4167f92d} /* (3, 21, 14) {real, imag} */,
  {32'hc199ab76, 32'h4276a5ca} /* (3, 21, 13) {real, imag} */,
  {32'h420ddc2a, 32'h41c51581} /* (3, 21, 12) {real, imag} */,
  {32'hc2b92c74, 32'h40071d10} /* (3, 21, 11) {real, imag} */,
  {32'h426ae4d5, 32'hc215a894} /* (3, 21, 10) {real, imag} */,
  {32'h42cb74d7, 32'h41b344a4} /* (3, 21, 9) {real, imag} */,
  {32'h3fa72650, 32'hc2939d9a} /* (3, 21, 8) {real, imag} */,
  {32'hc2c17232, 32'hc28f5583} /* (3, 21, 7) {real, imag} */,
  {32'hc20e735f, 32'hc28790fd} /* (3, 21, 6) {real, imag} */,
  {32'h4295ad7c, 32'h43003f30} /* (3, 21, 5) {real, imag} */,
  {32'h4263dc2e, 32'h42d23f48} /* (3, 21, 4) {real, imag} */,
  {32'hc281a59e, 32'h4247b68f} /* (3, 21, 3) {real, imag} */,
  {32'h43202238, 32'h42064858} /* (3, 21, 2) {real, imag} */,
  {32'hc3dbf8a2, 32'h432e74f4} /* (3, 21, 1) {real, imag} */,
  {32'h436a76db, 32'h00000000} /* (3, 21, 0) {real, imag} */,
  {32'h4425aeb0, 32'hc3aa32a8} /* (3, 20, 31) {real, imag} */,
  {32'hc3f4ea57, 32'hc190c25e} /* (3, 20, 30) {real, imag} */,
  {32'hc3720404, 32'h415bb653} /* (3, 20, 29) {real, imag} */,
  {32'h4328ef94, 32'hc2911b54} /* (3, 20, 28) {real, imag} */,
  {32'hc2eceb42, 32'hc319b204} /* (3, 20, 27) {real, imag} */,
  {32'hc083b4d4, 32'h4181253c} /* (3, 20, 26) {real, imag} */,
  {32'hc11ea0fa, 32'h42f45bcf} /* (3, 20, 25) {real, imag} */,
  {32'hc2b90d18, 32'h41a36a8f} /* (3, 20, 24) {real, imag} */,
  {32'h4298c029, 32'hc28f4550} /* (3, 20, 23) {real, imag} */,
  {32'h409f35aa, 32'h420c2f6b} /* (3, 20, 22) {real, imag} */,
  {32'hc321b0e4, 32'hbe2c1000} /* (3, 20, 21) {real, imag} */,
  {32'h41815652, 32'hc2ad4d62} /* (3, 20, 20) {real, imag} */,
  {32'h41f4c2db, 32'hc21bf312} /* (3, 20, 19) {real, imag} */,
  {32'h42527eaf, 32'h417a876a} /* (3, 20, 18) {real, imag} */,
  {32'h405b1db8, 32'hc0d526d6} /* (3, 20, 17) {real, imag} */,
  {32'hc325bce8, 32'h00000000} /* (3, 20, 16) {real, imag} */,
  {32'h405b1db8, 32'h40d526d6} /* (3, 20, 15) {real, imag} */,
  {32'h42527eaf, 32'hc17a876a} /* (3, 20, 14) {real, imag} */,
  {32'h41f4c2db, 32'h421bf312} /* (3, 20, 13) {real, imag} */,
  {32'h41815652, 32'h42ad4d62} /* (3, 20, 12) {real, imag} */,
  {32'hc321b0e4, 32'h3e2c1000} /* (3, 20, 11) {real, imag} */,
  {32'h409f35aa, 32'hc20c2f6b} /* (3, 20, 10) {real, imag} */,
  {32'h4298c029, 32'h428f4550} /* (3, 20, 9) {real, imag} */,
  {32'hc2b90d18, 32'hc1a36a8f} /* (3, 20, 8) {real, imag} */,
  {32'hc11ea0fa, 32'hc2f45bcf} /* (3, 20, 7) {real, imag} */,
  {32'hc083b4d4, 32'hc181253c} /* (3, 20, 6) {real, imag} */,
  {32'hc2eceb42, 32'h4319b204} /* (3, 20, 5) {real, imag} */,
  {32'h4328ef94, 32'h42911b54} /* (3, 20, 4) {real, imag} */,
  {32'hc3720404, 32'hc15bb653} /* (3, 20, 3) {real, imag} */,
  {32'hc3f4ea57, 32'h4190c25e} /* (3, 20, 2) {real, imag} */,
  {32'h4425aeb0, 32'h43aa32a8} /* (3, 20, 1) {real, imag} */,
  {32'h44730034, 32'h00000000} /* (3, 20, 0) {real, imag} */,
  {32'h449b8ef3, 32'hc398abfe} /* (3, 19, 31) {real, imag} */,
  {32'hc43aaa48, 32'h41c4d5d8} /* (3, 19, 30) {real, imag} */,
  {32'hc3461148, 32'h42058e1a} /* (3, 19, 29) {real, imag} */,
  {32'h438a32f5, 32'hc19f8964} /* (3, 19, 28) {real, imag} */,
  {32'hc31b8d9a, 32'h40f3d030} /* (3, 19, 27) {real, imag} */,
  {32'hc26c5ad8, 32'hc2682b13} /* (3, 19, 26) {real, imag} */,
  {32'h42f4c060, 32'h420c2202} /* (3, 19, 25) {real, imag} */,
  {32'hc1faa434, 32'h429a3efb} /* (3, 19, 24) {real, imag} */,
  {32'h42be1cd8, 32'hc11c547c} /* (3, 19, 23) {real, imag} */,
  {32'h41f817cc, 32'h415d98e0} /* (3, 19, 22) {real, imag} */,
  {32'hc35a0f76, 32'h4286f3fd} /* (3, 19, 21) {real, imag} */,
  {32'h40c339f8, 32'h40152ed0} /* (3, 19, 20) {real, imag} */,
  {32'h423242b5, 32'hc146fd80} /* (3, 19, 19) {real, imag} */,
  {32'h420da5f6, 32'h41ae7550} /* (3, 19, 18) {real, imag} */,
  {32'hc2436270, 32'hc1c0a79e} /* (3, 19, 17) {real, imag} */,
  {32'hc29b95a6, 32'h00000000} /* (3, 19, 16) {real, imag} */,
  {32'hc2436270, 32'h41c0a79e} /* (3, 19, 15) {real, imag} */,
  {32'h420da5f6, 32'hc1ae7550} /* (3, 19, 14) {real, imag} */,
  {32'h423242b5, 32'h4146fd80} /* (3, 19, 13) {real, imag} */,
  {32'h40c339f8, 32'hc0152ed0} /* (3, 19, 12) {real, imag} */,
  {32'hc35a0f76, 32'hc286f3fd} /* (3, 19, 11) {real, imag} */,
  {32'h41f817cc, 32'hc15d98e0} /* (3, 19, 10) {real, imag} */,
  {32'h42be1cd8, 32'h411c547c} /* (3, 19, 9) {real, imag} */,
  {32'hc1faa434, 32'hc29a3efb} /* (3, 19, 8) {real, imag} */,
  {32'h42f4c060, 32'hc20c2202} /* (3, 19, 7) {real, imag} */,
  {32'hc26c5ad8, 32'h42682b13} /* (3, 19, 6) {real, imag} */,
  {32'hc31b8d9a, 32'hc0f3d030} /* (3, 19, 5) {real, imag} */,
  {32'h438a32f5, 32'h419f8964} /* (3, 19, 4) {real, imag} */,
  {32'hc3461148, 32'hc2058e1a} /* (3, 19, 3) {real, imag} */,
  {32'hc43aaa48, 32'hc1c4d5d8} /* (3, 19, 2) {real, imag} */,
  {32'h449b8ef3, 32'h4398abfe} /* (3, 19, 1) {real, imag} */,
  {32'h44855cd5, 32'h00000000} /* (3, 19, 0) {real, imag} */,
  {32'h44c4da00, 32'hc3a64579} /* (3, 18, 31) {real, imag} */,
  {32'hc469b140, 32'h434edc60} /* (3, 18, 30) {real, imag} */,
  {32'hc343c27a, 32'hc1e91c1f} /* (3, 18, 29) {real, imag} */,
  {32'h4396c238, 32'hc2c6906c} /* (3, 18, 28) {real, imag} */,
  {32'hc33b046c, 32'h4314bbaf} /* (3, 18, 27) {real, imag} */,
  {32'hc2d827be, 32'hc24662e8} /* (3, 18, 26) {real, imag} */,
  {32'h41f6cd20, 32'hc18ccfa8} /* (3, 18, 25) {real, imag} */,
  {32'h4211e10a, 32'h421e859e} /* (3, 18, 24) {real, imag} */,
  {32'hc12085e2, 32'h4266fda2} /* (3, 18, 23) {real, imag} */,
  {32'h4281cd50, 32'hc26f1cee} /* (3, 18, 22) {real, imag} */,
  {32'hc2fbbd84, 32'h426fb701} /* (3, 18, 21) {real, imag} */,
  {32'h43297311, 32'hc299a3c7} /* (3, 18, 20) {real, imag} */,
  {32'hc31186b2, 32'hc27ad386} /* (3, 18, 19) {real, imag} */,
  {32'hc20285e7, 32'h43365e78} /* (3, 18, 18) {real, imag} */,
  {32'h41937f6b, 32'h41fa8c93} /* (3, 18, 17) {real, imag} */,
  {32'h429dcc5f, 32'h00000000} /* (3, 18, 16) {real, imag} */,
  {32'h41937f6b, 32'hc1fa8c93} /* (3, 18, 15) {real, imag} */,
  {32'hc20285e7, 32'hc3365e78} /* (3, 18, 14) {real, imag} */,
  {32'hc31186b2, 32'h427ad386} /* (3, 18, 13) {real, imag} */,
  {32'h43297311, 32'h4299a3c7} /* (3, 18, 12) {real, imag} */,
  {32'hc2fbbd84, 32'hc26fb701} /* (3, 18, 11) {real, imag} */,
  {32'h4281cd50, 32'h426f1cee} /* (3, 18, 10) {real, imag} */,
  {32'hc12085e2, 32'hc266fda2} /* (3, 18, 9) {real, imag} */,
  {32'h4211e10a, 32'hc21e859e} /* (3, 18, 8) {real, imag} */,
  {32'h41f6cd20, 32'h418ccfa8} /* (3, 18, 7) {real, imag} */,
  {32'hc2d827be, 32'h424662e8} /* (3, 18, 6) {real, imag} */,
  {32'hc33b046c, 32'hc314bbaf} /* (3, 18, 5) {real, imag} */,
  {32'h4396c238, 32'h42c6906c} /* (3, 18, 4) {real, imag} */,
  {32'hc343c27a, 32'h41e91c1f} /* (3, 18, 3) {real, imag} */,
  {32'hc469b140, 32'hc34edc60} /* (3, 18, 2) {real, imag} */,
  {32'h44c4da00, 32'h43a64579} /* (3, 18, 1) {real, imag} */,
  {32'h447a603a, 32'h00000000} /* (3, 18, 0) {real, imag} */,
  {32'h44d0ecee, 32'hc3895918} /* (3, 17, 31) {real, imag} */,
  {32'hc462778e, 32'h42b5f8ee} /* (3, 17, 30) {real, imag} */,
  {32'hc2d6ba25, 32'h41f7f168} /* (3, 17, 29) {real, imag} */,
  {32'h42bf8b10, 32'hc2c74668} /* (3, 17, 28) {real, imag} */,
  {32'hc2ebf0f0, 32'h407a4200} /* (3, 17, 27) {real, imag} */,
  {32'hc0574770, 32'hc2354137} /* (3, 17, 26) {real, imag} */,
  {32'h42c7569f, 32'hc3066c8a} /* (3, 17, 25) {real, imag} */,
  {32'hc234dd06, 32'h41f5fe40} /* (3, 17, 24) {real, imag} */,
  {32'h414c1714, 32'h42518e04} /* (3, 17, 23) {real, imag} */,
  {32'h4290b0b5, 32'hc1f48df5} /* (3, 17, 22) {real, imag} */,
  {32'hc1c3f7f4, 32'h42776145} /* (3, 17, 21) {real, imag} */,
  {32'hc26c4dee, 32'hc1cc4a9f} /* (3, 17, 20) {real, imag} */,
  {32'hc15476b0, 32'hc2650bbd} /* (3, 17, 19) {real, imag} */,
  {32'hc1cfe782, 32'h4273f2c9} /* (3, 17, 18) {real, imag} */,
  {32'h4259836d, 32'hc2180e0f} /* (3, 17, 17) {real, imag} */,
  {32'h41b4dd16, 32'h00000000} /* (3, 17, 16) {real, imag} */,
  {32'h4259836d, 32'h42180e0f} /* (3, 17, 15) {real, imag} */,
  {32'hc1cfe782, 32'hc273f2c9} /* (3, 17, 14) {real, imag} */,
  {32'hc15476b0, 32'h42650bbd} /* (3, 17, 13) {real, imag} */,
  {32'hc26c4dee, 32'h41cc4a9f} /* (3, 17, 12) {real, imag} */,
  {32'hc1c3f7f4, 32'hc2776145} /* (3, 17, 11) {real, imag} */,
  {32'h4290b0b5, 32'h41f48df5} /* (3, 17, 10) {real, imag} */,
  {32'h414c1714, 32'hc2518e04} /* (3, 17, 9) {real, imag} */,
  {32'hc234dd06, 32'hc1f5fe40} /* (3, 17, 8) {real, imag} */,
  {32'h42c7569f, 32'h43066c8a} /* (3, 17, 7) {real, imag} */,
  {32'hc0574770, 32'h42354137} /* (3, 17, 6) {real, imag} */,
  {32'hc2ebf0f0, 32'hc07a4200} /* (3, 17, 5) {real, imag} */,
  {32'h42bf8b10, 32'h42c74668} /* (3, 17, 4) {real, imag} */,
  {32'hc2d6ba25, 32'hc1f7f168} /* (3, 17, 3) {real, imag} */,
  {32'hc462778e, 32'hc2b5f8ee} /* (3, 17, 2) {real, imag} */,
  {32'h44d0ecee, 32'h43895918} /* (3, 17, 1) {real, imag} */,
  {32'h4484b9a4, 32'h00000000} /* (3, 17, 0) {real, imag} */,
  {32'h44ea1bb9, 32'hc359d10e} /* (3, 16, 31) {real, imag} */,
  {32'hc455d647, 32'h431bf9a8} /* (3, 16, 30) {real, imag} */,
  {32'h42fe41b8, 32'hc12884de} /* (3, 16, 29) {real, imag} */,
  {32'h4342840c, 32'hc2ab550b} /* (3, 16, 28) {real, imag} */,
  {32'hc320dd64, 32'h42952e7d} /* (3, 16, 27) {real, imag} */,
  {32'hc299ed7c, 32'hc2490adc} /* (3, 16, 26) {real, imag} */,
  {32'h41f24610, 32'hc22e9a62} /* (3, 16, 25) {real, imag} */,
  {32'hc2d7f3e6, 32'h42a9507a} /* (3, 16, 24) {real, imag} */,
  {32'h426be222, 32'h41f44ba4} /* (3, 16, 23) {real, imag} */,
  {32'hc22ed07c, 32'hc1930a55} /* (3, 16, 22) {real, imag} */,
  {32'h4115383c, 32'h428cf89c} /* (3, 16, 21) {real, imag} */,
  {32'hc1877651, 32'h42af3aba} /* (3, 16, 20) {real, imag} */,
  {32'h41b37304, 32'hc23e408c} /* (3, 16, 19) {real, imag} */,
  {32'h42d2a777, 32'h42a37ac5} /* (3, 16, 18) {real, imag} */,
  {32'hc177b108, 32'hc1aa5be3} /* (3, 16, 17) {real, imag} */,
  {32'h41faec94, 32'h00000000} /* (3, 16, 16) {real, imag} */,
  {32'hc177b108, 32'h41aa5be3} /* (3, 16, 15) {real, imag} */,
  {32'h42d2a777, 32'hc2a37ac5} /* (3, 16, 14) {real, imag} */,
  {32'h41b37304, 32'h423e408c} /* (3, 16, 13) {real, imag} */,
  {32'hc1877651, 32'hc2af3aba} /* (3, 16, 12) {real, imag} */,
  {32'h4115383c, 32'hc28cf89c} /* (3, 16, 11) {real, imag} */,
  {32'hc22ed07c, 32'h41930a55} /* (3, 16, 10) {real, imag} */,
  {32'h426be222, 32'hc1f44ba4} /* (3, 16, 9) {real, imag} */,
  {32'hc2d7f3e6, 32'hc2a9507a} /* (3, 16, 8) {real, imag} */,
  {32'h41f24610, 32'h422e9a62} /* (3, 16, 7) {real, imag} */,
  {32'hc299ed7c, 32'h42490adc} /* (3, 16, 6) {real, imag} */,
  {32'hc320dd64, 32'hc2952e7d} /* (3, 16, 5) {real, imag} */,
  {32'h4342840c, 32'h42ab550b} /* (3, 16, 4) {real, imag} */,
  {32'h42fe41b8, 32'h412884de} /* (3, 16, 3) {real, imag} */,
  {32'hc455d647, 32'hc31bf9a8} /* (3, 16, 2) {real, imag} */,
  {32'h44ea1bb9, 32'h4359d10e} /* (3, 16, 1) {real, imag} */,
  {32'h447db468, 32'h00000000} /* (3, 16, 0) {real, imag} */,
  {32'h44d42f2a, 32'hc3a494aa} /* (3, 15, 31) {real, imag} */,
  {32'hc44e0c26, 32'h435942d3} /* (3, 15, 30) {real, imag} */,
  {32'h42ad9605, 32'h419a2252} /* (3, 15, 29) {real, imag} */,
  {32'h4358386c, 32'hc2af05ee} /* (3, 15, 28) {real, imag} */,
  {32'hc34d9958, 32'h42bfa458} /* (3, 15, 27) {real, imag} */,
  {32'h42220c93, 32'hbf2d1d80} /* (3, 15, 26) {real, imag} */,
  {32'h426af63a, 32'hc2880f37} /* (3, 15, 25) {real, imag} */,
  {32'hc30f5e62, 32'h41910880} /* (3, 15, 24) {real, imag} */,
  {32'hc2181902, 32'hc06dd988} /* (3, 15, 23) {real, imag} */,
  {32'h41f4bfcc, 32'hc1d8019b} /* (3, 15, 22) {real, imag} */,
  {32'hc2756eea, 32'h41f24a76} /* (3, 15, 21) {real, imag} */,
  {32'h42927075, 32'hc1cc8e77} /* (3, 15, 20) {real, imag} */,
  {32'h428a14da, 32'hc165e3bc} /* (3, 15, 19) {real, imag} */,
  {32'h42ab91c6, 32'h3ef7e900} /* (3, 15, 18) {real, imag} */,
  {32'hc0f318f8, 32'h426ac249} /* (3, 15, 17) {real, imag} */,
  {32'hc2958154, 32'h00000000} /* (3, 15, 16) {real, imag} */,
  {32'hc0f318f8, 32'hc26ac249} /* (3, 15, 15) {real, imag} */,
  {32'h42ab91c6, 32'hbef7e900} /* (3, 15, 14) {real, imag} */,
  {32'h428a14da, 32'h4165e3bc} /* (3, 15, 13) {real, imag} */,
  {32'h42927075, 32'h41cc8e77} /* (3, 15, 12) {real, imag} */,
  {32'hc2756eea, 32'hc1f24a76} /* (3, 15, 11) {real, imag} */,
  {32'h41f4bfcc, 32'h41d8019b} /* (3, 15, 10) {real, imag} */,
  {32'hc2181902, 32'h406dd988} /* (3, 15, 9) {real, imag} */,
  {32'hc30f5e62, 32'hc1910880} /* (3, 15, 8) {real, imag} */,
  {32'h426af63a, 32'h42880f37} /* (3, 15, 7) {real, imag} */,
  {32'h42220c93, 32'h3f2d1d80} /* (3, 15, 6) {real, imag} */,
  {32'hc34d9958, 32'hc2bfa458} /* (3, 15, 5) {real, imag} */,
  {32'h4358386c, 32'h42af05ee} /* (3, 15, 4) {real, imag} */,
  {32'h42ad9605, 32'hc19a2252} /* (3, 15, 3) {real, imag} */,
  {32'hc44e0c26, 32'hc35942d3} /* (3, 15, 2) {real, imag} */,
  {32'h44d42f2a, 32'h43a494aa} /* (3, 15, 1) {real, imag} */,
  {32'h449c167a, 32'h00000000} /* (3, 15, 0) {real, imag} */,
  {32'h44d006fc, 32'hc3905243} /* (3, 14, 31) {real, imag} */,
  {32'hc453e808, 32'h42ee1bfb} /* (3, 14, 30) {real, imag} */,
  {32'h4341ff80, 32'h41c53c15} /* (3, 14, 29) {real, imag} */,
  {32'h4304389d, 32'hc32fdf5a} /* (3, 14, 28) {real, imag} */,
  {32'hc34fa836, 32'h438152a2} /* (3, 14, 27) {real, imag} */,
  {32'h42ac3332, 32'h4261967c} /* (3, 14, 26) {real, imag} */,
  {32'h42f367c8, 32'hc2da4bb3} /* (3, 14, 25) {real, imag} */,
  {32'hc2e2f24b, 32'h42a0a491} /* (3, 14, 24) {real, imag} */,
  {32'h41c102b5, 32'hc0e08e80} /* (3, 14, 23) {real, imag} */,
  {32'hc264065f, 32'h41a34800} /* (3, 14, 22) {real, imag} */,
  {32'h4231212c, 32'hc148081c} /* (3, 14, 21) {real, imag} */,
  {32'h4277b16c, 32'h4290994d} /* (3, 14, 20) {real, imag} */,
  {32'h410e5c50, 32'hc23c081a} /* (3, 14, 19) {real, imag} */,
  {32'hc213faf1, 32'h42aaf9e0} /* (3, 14, 18) {real, imag} */,
  {32'h428194d3, 32'hc222694a} /* (3, 14, 17) {real, imag} */,
  {32'h41982ffd, 32'h00000000} /* (3, 14, 16) {real, imag} */,
  {32'h428194d3, 32'h4222694a} /* (3, 14, 15) {real, imag} */,
  {32'hc213faf1, 32'hc2aaf9e0} /* (3, 14, 14) {real, imag} */,
  {32'h410e5c50, 32'h423c081a} /* (3, 14, 13) {real, imag} */,
  {32'h4277b16c, 32'hc290994d} /* (3, 14, 12) {real, imag} */,
  {32'h4231212c, 32'h4148081c} /* (3, 14, 11) {real, imag} */,
  {32'hc264065f, 32'hc1a34800} /* (3, 14, 10) {real, imag} */,
  {32'h41c102b5, 32'h40e08e80} /* (3, 14, 9) {real, imag} */,
  {32'hc2e2f24b, 32'hc2a0a491} /* (3, 14, 8) {real, imag} */,
  {32'h42f367c8, 32'h42da4bb3} /* (3, 14, 7) {real, imag} */,
  {32'h42ac3332, 32'hc261967c} /* (3, 14, 6) {real, imag} */,
  {32'hc34fa836, 32'hc38152a2} /* (3, 14, 5) {real, imag} */,
  {32'h4304389d, 32'h432fdf5a} /* (3, 14, 4) {real, imag} */,
  {32'h4341ff80, 32'hc1c53c15} /* (3, 14, 3) {real, imag} */,
  {32'hc453e808, 32'hc2ee1bfb} /* (3, 14, 2) {real, imag} */,
  {32'h44d006fc, 32'h43905243} /* (3, 14, 1) {real, imag} */,
  {32'h44a171b3, 32'h00000000} /* (3, 14, 0) {real, imag} */,
  {32'h44d33c3d, 32'hc3b15a3a} /* (3, 13, 31) {real, imag} */,
  {32'hc42fb5c0, 32'h420ad1ac} /* (3, 13, 30) {real, imag} */,
  {32'h43333b44, 32'h4121b558} /* (3, 13, 29) {real, imag} */,
  {32'h4336cd33, 32'hc31c777e} /* (3, 13, 28) {real, imag} */,
  {32'hc32cd4e4, 32'h432a7028} /* (3, 13, 27) {real, imag} */,
  {32'hc21d22fc, 32'h42f0f0c6} /* (3, 13, 26) {real, imag} */,
  {32'h41442830, 32'h428cd941} /* (3, 13, 25) {real, imag} */,
  {32'hc2def0fb, 32'h42e9c5fd} /* (3, 13, 24) {real, imag} */,
  {32'h42c82ac8, 32'h42cdd59e} /* (3, 13, 23) {real, imag} */,
  {32'hc2158f00, 32'hc230a39e} /* (3, 13, 22) {real, imag} */,
  {32'hc2106e82, 32'h42719352} /* (3, 13, 21) {real, imag} */,
  {32'hc2c7a176, 32'hc2d92b12} /* (3, 13, 20) {real, imag} */,
  {32'hc201362d, 32'h42fad6cc} /* (3, 13, 19) {real, imag} */,
  {32'h41569817, 32'h4202ed96} /* (3, 13, 18) {real, imag} */,
  {32'hc245b0c0, 32'h4296afce} /* (3, 13, 17) {real, imag} */,
  {32'hbea52c80, 32'h00000000} /* (3, 13, 16) {real, imag} */,
  {32'hc245b0c0, 32'hc296afce} /* (3, 13, 15) {real, imag} */,
  {32'h41569817, 32'hc202ed96} /* (3, 13, 14) {real, imag} */,
  {32'hc201362d, 32'hc2fad6cc} /* (3, 13, 13) {real, imag} */,
  {32'hc2c7a176, 32'h42d92b12} /* (3, 13, 12) {real, imag} */,
  {32'hc2106e82, 32'hc2719352} /* (3, 13, 11) {real, imag} */,
  {32'hc2158f00, 32'h4230a39e} /* (3, 13, 10) {real, imag} */,
  {32'h42c82ac8, 32'hc2cdd59e} /* (3, 13, 9) {real, imag} */,
  {32'hc2def0fb, 32'hc2e9c5fd} /* (3, 13, 8) {real, imag} */,
  {32'h41442830, 32'hc28cd941} /* (3, 13, 7) {real, imag} */,
  {32'hc21d22fc, 32'hc2f0f0c6} /* (3, 13, 6) {real, imag} */,
  {32'hc32cd4e4, 32'hc32a7028} /* (3, 13, 5) {real, imag} */,
  {32'h4336cd33, 32'h431c777e} /* (3, 13, 4) {real, imag} */,
  {32'h43333b44, 32'hc121b558} /* (3, 13, 3) {real, imag} */,
  {32'hc42fb5c0, 32'hc20ad1ac} /* (3, 13, 2) {real, imag} */,
  {32'h44d33c3d, 32'h43b15a3a} /* (3, 13, 1) {real, imag} */,
  {32'h44971ed1, 32'h00000000} /* (3, 13, 0) {real, imag} */,
  {32'h44b4d41c, 32'hc38021e4} /* (3, 12, 31) {real, imag} */,
  {32'hc4155e1a, 32'h41d75b1e} /* (3, 12, 30) {real, imag} */,
  {32'h43199eb6, 32'hc18bdcdf} /* (3, 12, 29) {real, imag} */,
  {32'h4312dea8, 32'hc2abaa9c} /* (3, 12, 28) {real, imag} */,
  {32'hc290b9ba, 32'h427215d2} /* (3, 12, 27) {real, imag} */,
  {32'hc237f14c, 32'h43425cae} /* (3, 12, 26) {real, imag} */,
  {32'hbf8e03b0, 32'h43023dd3} /* (3, 12, 25) {real, imag} */,
  {32'hc1ac1602, 32'h428c3670} /* (3, 12, 24) {real, imag} */,
  {32'h4265cbbe, 32'h427a8ddd} /* (3, 12, 23) {real, imag} */,
  {32'h4205439f, 32'hc0baaf52} /* (3, 12, 22) {real, imag} */,
  {32'hc2015ad0, 32'h430fd3be} /* (3, 12, 21) {real, imag} */,
  {32'hc1062771, 32'h4306326a} /* (3, 12, 20) {real, imag} */,
  {32'h4191c487, 32'hc18b802a} /* (3, 12, 19) {real, imag} */,
  {32'hc2db0f2a, 32'h428edd26} /* (3, 12, 18) {real, imag} */,
  {32'hc1ef1a75, 32'h413659bb} /* (3, 12, 17) {real, imag} */,
  {32'hc26feb98, 32'h00000000} /* (3, 12, 16) {real, imag} */,
  {32'hc1ef1a75, 32'hc13659bb} /* (3, 12, 15) {real, imag} */,
  {32'hc2db0f2a, 32'hc28edd26} /* (3, 12, 14) {real, imag} */,
  {32'h4191c487, 32'h418b802a} /* (3, 12, 13) {real, imag} */,
  {32'hc1062771, 32'hc306326a} /* (3, 12, 12) {real, imag} */,
  {32'hc2015ad0, 32'hc30fd3be} /* (3, 12, 11) {real, imag} */,
  {32'h4205439f, 32'h40baaf52} /* (3, 12, 10) {real, imag} */,
  {32'h4265cbbe, 32'hc27a8ddd} /* (3, 12, 9) {real, imag} */,
  {32'hc1ac1602, 32'hc28c3670} /* (3, 12, 8) {real, imag} */,
  {32'hbf8e03b0, 32'hc3023dd3} /* (3, 12, 7) {real, imag} */,
  {32'hc237f14c, 32'hc3425cae} /* (3, 12, 6) {real, imag} */,
  {32'hc290b9ba, 32'hc27215d2} /* (3, 12, 5) {real, imag} */,
  {32'h4312dea8, 32'h42abaa9c} /* (3, 12, 4) {real, imag} */,
  {32'h43199eb6, 32'h418bdcdf} /* (3, 12, 3) {real, imag} */,
  {32'hc4155e1a, 32'hc1d75b1e} /* (3, 12, 2) {real, imag} */,
  {32'h44b4d41c, 32'h438021e4} /* (3, 12, 1) {real, imag} */,
  {32'h4483458f, 32'h00000000} /* (3, 12, 0) {real, imag} */,
  {32'h4470b997, 32'hc220fb30} /* (3, 11, 31) {real, imag} */,
  {32'hc3ebb9be, 32'hc21db798} /* (3, 11, 30) {real, imag} */,
  {32'h425f7ead, 32'hc27f2aa7} /* (3, 11, 29) {real, imag} */,
  {32'h42ed4f3b, 32'hc2d07b2e} /* (3, 11, 28) {real, imag} */,
  {32'hc350046e, 32'h42d6b182} /* (3, 11, 27) {real, imag} */,
  {32'hc0c28b98, 32'h410967e8} /* (3, 11, 26) {real, imag} */,
  {32'h408482b8, 32'hc2a15d91} /* (3, 11, 25) {real, imag} */,
  {32'hc18ae4e3, 32'h42be47ac} /* (3, 11, 24) {real, imag} */,
  {32'h40cfc940, 32'hc2dc3447} /* (3, 11, 23) {real, imag} */,
  {32'hc23316e1, 32'h4297b37c} /* (3, 11, 22) {real, imag} */,
  {32'h424f7d31, 32'h42c81478} /* (3, 11, 21) {real, imag} */,
  {32'h41d5d553, 32'h4139285e} /* (3, 11, 20) {real, imag} */,
  {32'h41a2e35e, 32'hc21f1530} /* (3, 11, 19) {real, imag} */,
  {32'h40c1788e, 32'hc101e2ed} /* (3, 11, 18) {real, imag} */,
  {32'hc157a630, 32'h4181a5f8} /* (3, 11, 17) {real, imag} */,
  {32'h40aea346, 32'h00000000} /* (3, 11, 16) {real, imag} */,
  {32'hc157a630, 32'hc181a5f8} /* (3, 11, 15) {real, imag} */,
  {32'h40c1788e, 32'h4101e2ed} /* (3, 11, 14) {real, imag} */,
  {32'h41a2e35e, 32'h421f1530} /* (3, 11, 13) {real, imag} */,
  {32'h41d5d553, 32'hc139285e} /* (3, 11, 12) {real, imag} */,
  {32'h424f7d31, 32'hc2c81478} /* (3, 11, 11) {real, imag} */,
  {32'hc23316e1, 32'hc297b37c} /* (3, 11, 10) {real, imag} */,
  {32'h40cfc940, 32'h42dc3447} /* (3, 11, 9) {real, imag} */,
  {32'hc18ae4e3, 32'hc2be47ac} /* (3, 11, 8) {real, imag} */,
  {32'h408482b8, 32'h42a15d91} /* (3, 11, 7) {real, imag} */,
  {32'hc0c28b98, 32'hc10967e8} /* (3, 11, 6) {real, imag} */,
  {32'hc350046e, 32'hc2d6b182} /* (3, 11, 5) {real, imag} */,
  {32'h42ed4f3b, 32'h42d07b2e} /* (3, 11, 4) {real, imag} */,
  {32'h425f7ead, 32'h427f2aa7} /* (3, 11, 3) {real, imag} */,
  {32'hc3ebb9be, 32'h421db798} /* (3, 11, 2) {real, imag} */,
  {32'h4470b997, 32'h4220fb30} /* (3, 11, 1) {real, imag} */,
  {32'h441f28c5, 32'h00000000} /* (3, 11, 0) {real, imag} */,
  {32'hc32fba58, 32'h4294f587} /* (3, 10, 31) {real, imag} */,
  {32'h42c2f5c0, 32'hc2ec1e7a} /* (3, 10, 30) {real, imag} */,
  {32'h42032eee, 32'hc3335521} /* (3, 10, 29) {real, imag} */,
  {32'hc17e7d54, 32'h42296a96} /* (3, 10, 28) {real, imag} */,
  {32'hc1fae384, 32'hc219e607} /* (3, 10, 27) {real, imag} */,
  {32'h42ab4608, 32'h420cca80} /* (3, 10, 26) {real, imag} */,
  {32'hc23ecb82, 32'h41f58c8e} /* (3, 10, 25) {real, imag} */,
  {32'h416f1c56, 32'h41da35d6} /* (3, 10, 24) {real, imag} */,
  {32'h41d57a02, 32'h3f25fc00} /* (3, 10, 23) {real, imag} */,
  {32'h3fb93d80, 32'h41a57f18} /* (3, 10, 22) {real, imag} */,
  {32'hc291aa80, 32'hc1eaf942} /* (3, 10, 21) {real, imag} */,
  {32'hc276135e, 32'h40dc31c0} /* (3, 10, 20) {real, imag} */,
  {32'hc283e88c, 32'h42254c40} /* (3, 10, 19) {real, imag} */,
  {32'h42da4813, 32'hc25eee68} /* (3, 10, 18) {real, imag} */,
  {32'hc2bfc774, 32'hc25a6675} /* (3, 10, 17) {real, imag} */,
  {32'hc238b40d, 32'h00000000} /* (3, 10, 16) {real, imag} */,
  {32'hc2bfc774, 32'h425a6675} /* (3, 10, 15) {real, imag} */,
  {32'h42da4813, 32'h425eee68} /* (3, 10, 14) {real, imag} */,
  {32'hc283e88c, 32'hc2254c40} /* (3, 10, 13) {real, imag} */,
  {32'hc276135e, 32'hc0dc31c0} /* (3, 10, 12) {real, imag} */,
  {32'hc291aa80, 32'h41eaf942} /* (3, 10, 11) {real, imag} */,
  {32'h3fb93d80, 32'hc1a57f18} /* (3, 10, 10) {real, imag} */,
  {32'h41d57a02, 32'hbf25fc00} /* (3, 10, 9) {real, imag} */,
  {32'h416f1c56, 32'hc1da35d6} /* (3, 10, 8) {real, imag} */,
  {32'hc23ecb82, 32'hc1f58c8e} /* (3, 10, 7) {real, imag} */,
  {32'h42ab4608, 32'hc20cca80} /* (3, 10, 6) {real, imag} */,
  {32'hc1fae384, 32'h4219e607} /* (3, 10, 5) {real, imag} */,
  {32'hc17e7d54, 32'hc2296a96} /* (3, 10, 4) {real, imag} */,
  {32'h42032eee, 32'h43335521} /* (3, 10, 3) {real, imag} */,
  {32'h42c2f5c0, 32'h42ec1e7a} /* (3, 10, 2) {real, imag} */,
  {32'hc32fba58, 32'hc294f587} /* (3, 10, 1) {real, imag} */,
  {32'hc2c69c54, 32'h00000000} /* (3, 10, 0) {real, imag} */,
  {32'hc475d5df, 32'h42c76e2d} /* (3, 9, 31) {real, imag} */,
  {32'h43e5e7b2, 32'hc35d8e1c} /* (3, 9, 30) {real, imag} */,
  {32'h41f7f520, 32'hc2245e08} /* (3, 9, 29) {real, imag} */,
  {32'hc258a7e4, 32'h42c3e883} /* (3, 9, 28) {real, imag} */,
  {32'h43421ec0, 32'hc3204236} /* (3, 9, 27) {real, imag} */,
  {32'h425aefe3, 32'h42d06ba9} /* (3, 9, 26) {real, imag} */,
  {32'hc2d45b86, 32'h42214f88} /* (3, 9, 25) {real, imag} */,
  {32'h4308bc84, 32'hc22ef991} /* (3, 9, 24) {real, imag} */,
  {32'h42522a24, 32'h419ab55f} /* (3, 9, 23) {real, imag} */,
  {32'hc24a82c4, 32'hc20f996e} /* (3, 9, 22) {real, imag} */,
  {32'h41b86ae1, 32'hc22f38a9} /* (3, 9, 21) {real, imag} */,
  {32'hc1d0f1ed, 32'hc168878c} /* (3, 9, 20) {real, imag} */,
  {32'h425ea9d6, 32'hc328a150} /* (3, 9, 19) {real, imag} */,
  {32'h427e6312, 32'h42852a1e} /* (3, 9, 18) {real, imag} */,
  {32'hc21a74b2, 32'hc25e79ca} /* (3, 9, 17) {real, imag} */,
  {32'hc186f04b, 32'h00000000} /* (3, 9, 16) {real, imag} */,
  {32'hc21a74b2, 32'h425e79ca} /* (3, 9, 15) {real, imag} */,
  {32'h427e6312, 32'hc2852a1e} /* (3, 9, 14) {real, imag} */,
  {32'h425ea9d6, 32'h4328a150} /* (3, 9, 13) {real, imag} */,
  {32'hc1d0f1ed, 32'h4168878c} /* (3, 9, 12) {real, imag} */,
  {32'h41b86ae1, 32'h422f38a9} /* (3, 9, 11) {real, imag} */,
  {32'hc24a82c4, 32'h420f996e} /* (3, 9, 10) {real, imag} */,
  {32'h42522a24, 32'hc19ab55f} /* (3, 9, 9) {real, imag} */,
  {32'h4308bc84, 32'h422ef991} /* (3, 9, 8) {real, imag} */,
  {32'hc2d45b86, 32'hc2214f88} /* (3, 9, 7) {real, imag} */,
  {32'h425aefe3, 32'hc2d06ba9} /* (3, 9, 6) {real, imag} */,
  {32'h43421ec0, 32'h43204236} /* (3, 9, 5) {real, imag} */,
  {32'hc258a7e4, 32'hc2c3e883} /* (3, 9, 4) {real, imag} */,
  {32'h41f7f520, 32'h42245e08} /* (3, 9, 3) {real, imag} */,
  {32'h43e5e7b2, 32'h435d8e1c} /* (3, 9, 2) {real, imag} */,
  {32'hc475d5df, 32'hc2c76e2d} /* (3, 9, 1) {real, imag} */,
  {32'hc3d6a2ac, 32'h00000000} /* (3, 9, 0) {real, imag} */,
  {32'hc4995621, 32'h41ca1510} /* (3, 8, 31) {real, imag} */,
  {32'h4431c39e, 32'hc110d4c4} /* (3, 8, 30) {real, imag} */,
  {32'h42cc96c7, 32'hc2206622} /* (3, 8, 29) {real, imag} */,
  {32'hc30d4696, 32'hc29f0de0} /* (3, 8, 28) {real, imag} */,
  {32'h4360835d, 32'hc31d1722} /* (3, 8, 27) {real, imag} */,
  {32'hc19e44e5, 32'h428d1c3c} /* (3, 8, 26) {real, imag} */,
  {32'hc29a713a, 32'h420cd578} /* (3, 8, 25) {real, imag} */,
  {32'h42533db4, 32'hc2b5540c} /* (3, 8, 24) {real, imag} */,
  {32'h425b1c4c, 32'h42f78c47} /* (3, 8, 23) {real, imag} */,
  {32'hc2c3308c, 32'hc317ec0a} /* (3, 8, 22) {real, imag} */,
  {32'h4214e5aa, 32'h4242c243} /* (3, 8, 21) {real, imag} */,
  {32'hc2a82682, 32'hc194ea9d} /* (3, 8, 20) {real, imag} */,
  {32'h420871ca, 32'hc2b912fd} /* (3, 8, 19) {real, imag} */,
  {32'h423ec7dd, 32'hc1c18933} /* (3, 8, 18) {real, imag} */,
  {32'h41b5fe58, 32'h418b3c50} /* (3, 8, 17) {real, imag} */,
  {32'hc1672c67, 32'h00000000} /* (3, 8, 16) {real, imag} */,
  {32'h41b5fe58, 32'hc18b3c50} /* (3, 8, 15) {real, imag} */,
  {32'h423ec7dd, 32'h41c18933} /* (3, 8, 14) {real, imag} */,
  {32'h420871ca, 32'h42b912fd} /* (3, 8, 13) {real, imag} */,
  {32'hc2a82682, 32'h4194ea9d} /* (3, 8, 12) {real, imag} */,
  {32'h4214e5aa, 32'hc242c243} /* (3, 8, 11) {real, imag} */,
  {32'hc2c3308c, 32'h4317ec0a} /* (3, 8, 10) {real, imag} */,
  {32'h425b1c4c, 32'hc2f78c47} /* (3, 8, 9) {real, imag} */,
  {32'h42533db4, 32'h42b5540c} /* (3, 8, 8) {real, imag} */,
  {32'hc29a713a, 32'hc20cd578} /* (3, 8, 7) {real, imag} */,
  {32'hc19e44e5, 32'hc28d1c3c} /* (3, 8, 6) {real, imag} */,
  {32'h4360835d, 32'h431d1722} /* (3, 8, 5) {real, imag} */,
  {32'hc30d4696, 32'h429f0de0} /* (3, 8, 4) {real, imag} */,
  {32'h42cc96c7, 32'h42206622} /* (3, 8, 3) {real, imag} */,
  {32'h4431c39e, 32'h4110d4c4} /* (3, 8, 2) {real, imag} */,
  {32'hc4995621, 32'hc1ca1510} /* (3, 8, 1) {real, imag} */,
  {32'hc42f3e6f, 32'h00000000} /* (3, 8, 0) {real, imag} */,
  {32'hc4aeb2e6, 32'h437c74f6} /* (3, 7, 31) {real, imag} */,
  {32'h44410b06, 32'h42927bc8} /* (3, 7, 30) {real, imag} */,
  {32'h432836b1, 32'hc29dff4f} /* (3, 7, 29) {real, imag} */,
  {32'h42426298, 32'hc3133b96} /* (3, 7, 28) {real, imag} */,
  {32'h435081d4, 32'hc3282ec3} /* (3, 7, 27) {real, imag} */,
  {32'h41834a6a, 32'h42c49e7c} /* (3, 7, 26) {real, imag} */,
  {32'hc2d7bfc0, 32'h41cd160e} /* (3, 7, 25) {real, imag} */,
  {32'h421317ac, 32'h42256ca2} /* (3, 7, 24) {real, imag} */,
  {32'hc2021d21, 32'h4117b11f} /* (3, 7, 23) {real, imag} */,
  {32'hc2c08a51, 32'h428db4b6} /* (3, 7, 22) {real, imag} */,
  {32'hc192ffd8, 32'hc28bafb4} /* (3, 7, 21) {real, imag} */,
  {32'h408cbbc4, 32'h430cfa75} /* (3, 7, 20) {real, imag} */,
  {32'h4274f530, 32'hc24228c7} /* (3, 7, 19) {real, imag} */,
  {32'h40dab9c2, 32'hc29dfd2a} /* (3, 7, 18) {real, imag} */,
  {32'hbff2f600, 32'hc2fd5354} /* (3, 7, 17) {real, imag} */,
  {32'h4289b344, 32'h00000000} /* (3, 7, 16) {real, imag} */,
  {32'hbff2f600, 32'h42fd5354} /* (3, 7, 15) {real, imag} */,
  {32'h40dab9c2, 32'h429dfd2a} /* (3, 7, 14) {real, imag} */,
  {32'h4274f530, 32'h424228c7} /* (3, 7, 13) {real, imag} */,
  {32'h408cbbc4, 32'hc30cfa75} /* (3, 7, 12) {real, imag} */,
  {32'hc192ffd8, 32'h428bafb4} /* (3, 7, 11) {real, imag} */,
  {32'hc2c08a51, 32'hc28db4b6} /* (3, 7, 10) {real, imag} */,
  {32'hc2021d21, 32'hc117b11f} /* (3, 7, 9) {real, imag} */,
  {32'h421317ac, 32'hc2256ca2} /* (3, 7, 8) {real, imag} */,
  {32'hc2d7bfc0, 32'hc1cd160e} /* (3, 7, 7) {real, imag} */,
  {32'h41834a6a, 32'hc2c49e7c} /* (3, 7, 6) {real, imag} */,
  {32'h435081d4, 32'h43282ec3} /* (3, 7, 5) {real, imag} */,
  {32'h42426298, 32'h43133b96} /* (3, 7, 4) {real, imag} */,
  {32'h432836b1, 32'h429dff4f} /* (3, 7, 3) {real, imag} */,
  {32'h44410b06, 32'hc2927bc8} /* (3, 7, 2) {real, imag} */,
  {32'hc4aeb2e6, 32'hc37c74f6} /* (3, 7, 1) {real, imag} */,
  {32'hc43a6d5d, 32'h00000000} /* (3, 7, 0) {real, imag} */,
  {32'hc4a15e22, 32'h440520fa} /* (3, 6, 31) {real, imag} */,
  {32'h4405a61e, 32'hc283072e} /* (3, 6, 30) {real, imag} */,
  {32'h4336d7d4, 32'hc24769ea} /* (3, 6, 29) {real, imag} */,
  {32'hc2110544, 32'hc3226951} /* (3, 6, 28) {real, imag} */,
  {32'h42937296, 32'hc25b8e63} /* (3, 6, 27) {real, imag} */,
  {32'h40008430, 32'hc29ef5e4} /* (3, 6, 26) {real, imag} */,
  {32'hc11d9e38, 32'hc27e31ff} /* (3, 6, 25) {real, imag} */,
  {32'h42db9e08, 32'hc2d3e76a} /* (3, 6, 24) {real, imag} */,
  {32'h42e2f856, 32'h4226aaf4} /* (3, 6, 23) {real, imag} */,
  {32'hc2413639, 32'h4269ec25} /* (3, 6, 22) {real, imag} */,
  {32'h41e1ffbe, 32'hc2b87a0c} /* (3, 6, 21) {real, imag} */,
  {32'h3fa4a0c0, 32'h41b8fead} /* (3, 6, 20) {real, imag} */,
  {32'hc27dc770, 32'hc1f35578} /* (3, 6, 19) {real, imag} */,
  {32'hc0abc25c, 32'hc07e72f8} /* (3, 6, 18) {real, imag} */,
  {32'h410499dc, 32'h4280a599} /* (3, 6, 17) {real, imag} */,
  {32'hc26d5ffc, 32'h00000000} /* (3, 6, 16) {real, imag} */,
  {32'h410499dc, 32'hc280a599} /* (3, 6, 15) {real, imag} */,
  {32'hc0abc25c, 32'h407e72f8} /* (3, 6, 14) {real, imag} */,
  {32'hc27dc770, 32'h41f35578} /* (3, 6, 13) {real, imag} */,
  {32'h3fa4a0c0, 32'hc1b8fead} /* (3, 6, 12) {real, imag} */,
  {32'h41e1ffbe, 32'h42b87a0c} /* (3, 6, 11) {real, imag} */,
  {32'hc2413639, 32'hc269ec25} /* (3, 6, 10) {real, imag} */,
  {32'h42e2f856, 32'hc226aaf4} /* (3, 6, 9) {real, imag} */,
  {32'h42db9e08, 32'h42d3e76a} /* (3, 6, 8) {real, imag} */,
  {32'hc11d9e38, 32'h427e31ff} /* (3, 6, 7) {real, imag} */,
  {32'h40008430, 32'h429ef5e4} /* (3, 6, 6) {real, imag} */,
  {32'h42937296, 32'h425b8e63} /* (3, 6, 5) {real, imag} */,
  {32'hc2110544, 32'h43226951} /* (3, 6, 4) {real, imag} */,
  {32'h4336d7d4, 32'h424769ea} /* (3, 6, 3) {real, imag} */,
  {32'h4405a61e, 32'h4283072e} /* (3, 6, 2) {real, imag} */,
  {32'hc4a15e22, 32'hc40520fa} /* (3, 6, 1) {real, imag} */,
  {32'hc42a6f7a, 32'h00000000} /* (3, 6, 0) {real, imag} */,
  {32'hc47734e0, 32'h448125c0} /* (3, 5, 31) {real, imag} */,
  {32'h431f3532, 32'hc34fba76} /* (3, 5, 30) {real, imag} */,
  {32'h4396c1cb, 32'hc1c28af8} /* (3, 5, 29) {real, imag} */,
  {32'hc2b4db3b, 32'hc31e978b} /* (3, 5, 28) {real, imag} */,
  {32'h42800f75, 32'h413b97b8} /* (3, 5, 27) {real, imag} */,
  {32'h429f156f, 32'h41a0b5b8} /* (3, 5, 26) {real, imag} */,
  {32'h4259213a, 32'hc21549ea} /* (3, 5, 25) {real, imag} */,
  {32'hc29ec2d6, 32'hc284983c} /* (3, 5, 24) {real, imag} */,
  {32'h422c074e, 32'h41c9d869} /* (3, 5, 23) {real, imag} */,
  {32'h42808f5a, 32'h3d8a0200} /* (3, 5, 22) {real, imag} */,
  {32'hc2a3fe6c, 32'h419b48a7} /* (3, 5, 21) {real, imag} */,
  {32'hc0f1ab70, 32'hc26dff78} /* (3, 5, 20) {real, imag} */,
  {32'h41c589ba, 32'h41c84fa2} /* (3, 5, 19) {real, imag} */,
  {32'h4114be8a, 32'h429ca830} /* (3, 5, 18) {real, imag} */,
  {32'hc23a89e4, 32'hc281ed82} /* (3, 5, 17) {real, imag} */,
  {32'hc122d85a, 32'h00000000} /* (3, 5, 16) {real, imag} */,
  {32'hc23a89e4, 32'h4281ed82} /* (3, 5, 15) {real, imag} */,
  {32'h4114be8a, 32'hc29ca830} /* (3, 5, 14) {real, imag} */,
  {32'h41c589ba, 32'hc1c84fa2} /* (3, 5, 13) {real, imag} */,
  {32'hc0f1ab70, 32'h426dff78} /* (3, 5, 12) {real, imag} */,
  {32'hc2a3fe6c, 32'hc19b48a7} /* (3, 5, 11) {real, imag} */,
  {32'h42808f5a, 32'hbd8a0200} /* (3, 5, 10) {real, imag} */,
  {32'h422c074e, 32'hc1c9d869} /* (3, 5, 9) {real, imag} */,
  {32'hc29ec2d6, 32'h4284983c} /* (3, 5, 8) {real, imag} */,
  {32'h4259213a, 32'h421549ea} /* (3, 5, 7) {real, imag} */,
  {32'h429f156f, 32'hc1a0b5b8} /* (3, 5, 6) {real, imag} */,
  {32'h42800f75, 32'hc13b97b8} /* (3, 5, 5) {real, imag} */,
  {32'hc2b4db3b, 32'h431e978b} /* (3, 5, 4) {real, imag} */,
  {32'h4396c1cb, 32'h41c28af8} /* (3, 5, 3) {real, imag} */,
  {32'h431f3532, 32'h434fba76} /* (3, 5, 2) {real, imag} */,
  {32'hc47734e0, 32'hc48125c0} /* (3, 5, 1) {real, imag} */,
  {32'hc405f6b8, 32'h00000000} /* (3, 5, 0) {real, imag} */,
  {32'hc4523ef2, 32'h44baa9e8} /* (3, 4, 31) {real, imag} */,
  {32'hc322463e, 32'hc37e736c} /* (3, 4, 30) {real, imag} */,
  {32'h436255ad, 32'h42a4e42c} /* (3, 4, 29) {real, imag} */,
  {32'h4280c424, 32'hc36c638a} /* (3, 4, 28) {real, imag} */,
  {32'h4317c1f3, 32'h426e53d2} /* (3, 4, 27) {real, imag} */,
  {32'h42718f9c, 32'hc1cb57c6} /* (3, 4, 26) {real, imag} */,
  {32'hc2276aa4, 32'h41bd74e8} /* (3, 4, 25) {real, imag} */,
  {32'h4150aa34, 32'h4266762c} /* (3, 4, 24) {real, imag} */,
  {32'h4247bd53, 32'hc24ccbb5} /* (3, 4, 23) {real, imag} */,
  {32'h40f1cf50, 32'hc27cea61} /* (3, 4, 22) {real, imag} */,
  {32'h41ac0dd4, 32'h42907a73} /* (3, 4, 21) {real, imag} */,
  {32'h4223f8fb, 32'hc24236fc} /* (3, 4, 20) {real, imag} */,
  {32'h41b4b4e7, 32'h424905f0} /* (3, 4, 19) {real, imag} */,
  {32'hc14e43f4, 32'hc1a85a62} /* (3, 4, 18) {real, imag} */,
  {32'h414617e0, 32'hc1ec38a4} /* (3, 4, 17) {real, imag} */,
  {32'h42965d82, 32'h00000000} /* (3, 4, 16) {real, imag} */,
  {32'h414617e0, 32'h41ec38a4} /* (3, 4, 15) {real, imag} */,
  {32'hc14e43f4, 32'h41a85a62} /* (3, 4, 14) {real, imag} */,
  {32'h41b4b4e7, 32'hc24905f0} /* (3, 4, 13) {real, imag} */,
  {32'h4223f8fb, 32'h424236fc} /* (3, 4, 12) {real, imag} */,
  {32'h41ac0dd4, 32'hc2907a73} /* (3, 4, 11) {real, imag} */,
  {32'h40f1cf50, 32'h427cea61} /* (3, 4, 10) {real, imag} */,
  {32'h4247bd53, 32'h424ccbb5} /* (3, 4, 9) {real, imag} */,
  {32'h4150aa34, 32'hc266762c} /* (3, 4, 8) {real, imag} */,
  {32'hc2276aa4, 32'hc1bd74e8} /* (3, 4, 7) {real, imag} */,
  {32'h42718f9c, 32'h41cb57c6} /* (3, 4, 6) {real, imag} */,
  {32'h4317c1f3, 32'hc26e53d2} /* (3, 4, 5) {real, imag} */,
  {32'h4280c424, 32'h436c638a} /* (3, 4, 4) {real, imag} */,
  {32'h436255ad, 32'hc2a4e42c} /* (3, 4, 3) {real, imag} */,
  {32'hc322463e, 32'h437e736c} /* (3, 4, 2) {real, imag} */,
  {32'hc4523ef2, 32'hc4baa9e8} /* (3, 4, 1) {real, imag} */,
  {32'hc3b805ed, 32'h00000000} /* (3, 4, 0) {real, imag} */,
  {32'hc436cc18, 32'h44c10ebc} /* (3, 3, 31) {real, imag} */,
  {32'hc3ae1108, 32'hc3eda99b} /* (3, 3, 30) {real, imag} */,
  {32'h436b30aa, 32'h429ed403} /* (3, 3, 29) {real, imag} */,
  {32'h421af264, 32'hc35cb320} /* (3, 3, 28) {real, imag} */,
  {32'h435cd293, 32'h4221f893} /* (3, 3, 27) {real, imag} */,
  {32'h42a3cd7d, 32'hc15e6610} /* (3, 3, 26) {real, imag} */,
  {32'h428d7a84, 32'hc1e70430} /* (3, 3, 25) {real, imag} */,
  {32'hc1de8c02, 32'hc270b10c} /* (3, 3, 24) {real, imag} */,
  {32'h41070e1c, 32'hc28ddd42} /* (3, 3, 23) {real, imag} */,
  {32'hc09bef9c, 32'hc296b52d} /* (3, 3, 22) {real, imag} */,
  {32'h3e709b00, 32'hc227c3bc} /* (3, 3, 21) {real, imag} */,
  {32'hc2391efc, 32'hc221955c} /* (3, 3, 20) {real, imag} */,
  {32'h42172b29, 32'h416c6c10} /* (3, 3, 19) {real, imag} */,
  {32'hc285cbc8, 32'h419f947c} /* (3, 3, 18) {real, imag} */,
  {32'h42c20db1, 32'hc2980ee2} /* (3, 3, 17) {real, imag} */,
  {32'h42410bf4, 32'h00000000} /* (3, 3, 16) {real, imag} */,
  {32'h42c20db1, 32'h42980ee2} /* (3, 3, 15) {real, imag} */,
  {32'hc285cbc8, 32'hc19f947c} /* (3, 3, 14) {real, imag} */,
  {32'h42172b29, 32'hc16c6c10} /* (3, 3, 13) {real, imag} */,
  {32'hc2391efc, 32'h4221955c} /* (3, 3, 12) {real, imag} */,
  {32'h3e709b00, 32'h4227c3bc} /* (3, 3, 11) {real, imag} */,
  {32'hc09bef9c, 32'h4296b52d} /* (3, 3, 10) {real, imag} */,
  {32'h41070e1c, 32'h428ddd42} /* (3, 3, 9) {real, imag} */,
  {32'hc1de8c02, 32'h4270b10c} /* (3, 3, 8) {real, imag} */,
  {32'h428d7a84, 32'h41e70430} /* (3, 3, 7) {real, imag} */,
  {32'h42a3cd7d, 32'h415e6610} /* (3, 3, 6) {real, imag} */,
  {32'h435cd293, 32'hc221f893} /* (3, 3, 5) {real, imag} */,
  {32'h421af264, 32'h435cb320} /* (3, 3, 4) {real, imag} */,
  {32'h436b30aa, 32'hc29ed403} /* (3, 3, 3) {real, imag} */,
  {32'hc3ae1108, 32'h43eda99b} /* (3, 3, 2) {real, imag} */,
  {32'hc436cc18, 32'hc4c10ebc} /* (3, 3, 1) {real, imag} */,
  {32'hc3f6eb4c, 32'h00000000} /* (3, 3, 0) {real, imag} */,
  {32'hc416e6cf, 32'h44b2dbca} /* (3, 2, 31) {real, imag} */,
  {32'hc3b87d18, 32'hc4086084} /* (3, 2, 30) {real, imag} */,
  {32'h4324d781, 32'h42ec0f21} /* (3, 2, 29) {real, imag} */,
  {32'h432894c0, 32'hc3628f22} /* (3, 2, 28) {real, imag} */,
  {32'h42a9adb9, 32'h4292e8c4} /* (3, 2, 27) {real, imag} */,
  {32'h42cb4088, 32'h4190210e} /* (3, 2, 26) {real, imag} */,
  {32'h42976e7e, 32'h429dae5a} /* (3, 2, 25) {real, imag} */,
  {32'hc2e8b24f, 32'hc2946677} /* (3, 2, 24) {real, imag} */,
  {32'h42008ea2, 32'hc29caff0} /* (3, 2, 23) {real, imag} */,
  {32'h41fa6feb, 32'hc2490322} /* (3, 2, 22) {real, imag} */,
  {32'h42b5e5a5, 32'h421b70b1} /* (3, 2, 21) {real, imag} */,
  {32'h405b23e8, 32'h4258a1ae} /* (3, 2, 20) {real, imag} */,
  {32'hc2b8c8f9, 32'hc1ee55af} /* (3, 2, 19) {real, imag} */,
  {32'h40740774, 32'h427b6ac5} /* (3, 2, 18) {real, imag} */,
  {32'hc18b2626, 32'h41d1ab0c} /* (3, 2, 17) {real, imag} */,
  {32'hbe7dd180, 32'h00000000} /* (3, 2, 16) {real, imag} */,
  {32'hc18b2626, 32'hc1d1ab0c} /* (3, 2, 15) {real, imag} */,
  {32'h40740774, 32'hc27b6ac5} /* (3, 2, 14) {real, imag} */,
  {32'hc2b8c8f9, 32'h41ee55af} /* (3, 2, 13) {real, imag} */,
  {32'h405b23e8, 32'hc258a1ae} /* (3, 2, 12) {real, imag} */,
  {32'h42b5e5a5, 32'hc21b70b1} /* (3, 2, 11) {real, imag} */,
  {32'h41fa6feb, 32'h42490322} /* (3, 2, 10) {real, imag} */,
  {32'h42008ea2, 32'h429caff0} /* (3, 2, 9) {real, imag} */,
  {32'hc2e8b24f, 32'h42946677} /* (3, 2, 8) {real, imag} */,
  {32'h42976e7e, 32'hc29dae5a} /* (3, 2, 7) {real, imag} */,
  {32'h42cb4088, 32'hc190210e} /* (3, 2, 6) {real, imag} */,
  {32'h42a9adb9, 32'hc292e8c4} /* (3, 2, 5) {real, imag} */,
  {32'h432894c0, 32'h43628f22} /* (3, 2, 4) {real, imag} */,
  {32'h4324d781, 32'hc2ec0f21} /* (3, 2, 3) {real, imag} */,
  {32'hc3b87d18, 32'h44086084} /* (3, 2, 2) {real, imag} */,
  {32'hc416e6cf, 32'hc4b2dbca} /* (3, 2, 1) {real, imag} */,
  {32'hc37883b6, 32'h00000000} /* (3, 2, 0) {real, imag} */,
  {32'hc41281ab, 32'h44a143f0} /* (3, 1, 31) {real, imag} */,
  {32'hc3b2aa4d, 32'hc3fd2d6b} /* (3, 1, 30) {real, imag} */,
  {32'h429dfe6a, 32'hc205c217} /* (3, 1, 29) {real, imag} */,
  {32'h42ec2c6b, 32'hc38620c7} /* (3, 1, 28) {real, imag} */,
  {32'h43019672, 32'hc29fca6f} /* (3, 1, 27) {real, imag} */,
  {32'h41cae78c, 32'h42a5c8b8} /* (3, 1, 26) {real, imag} */,
  {32'h41ac97fc, 32'h4289026a} /* (3, 1, 25) {real, imag} */,
  {32'hc29d4c87, 32'hc3118d27} /* (3, 1, 24) {real, imag} */,
  {32'h4200fe80, 32'hc2d32d16} /* (3, 1, 23) {real, imag} */,
  {32'h429e5cff, 32'hc1d4dd10} /* (3, 1, 22) {real, imag} */,
  {32'h416275d2, 32'hc1ca126e} /* (3, 1, 21) {real, imag} */,
  {32'hc24ca7c8, 32'hc236d2aa} /* (3, 1, 20) {real, imag} */,
  {32'h423e5143, 32'h41389732} /* (3, 1, 19) {real, imag} */,
  {32'hc1cf5cf6, 32'hc17e4bb8} /* (3, 1, 18) {real, imag} */,
  {32'h42276aeb, 32'h40bba264} /* (3, 1, 17) {real, imag} */,
  {32'h425ff871, 32'h00000000} /* (3, 1, 16) {real, imag} */,
  {32'h42276aeb, 32'hc0bba264} /* (3, 1, 15) {real, imag} */,
  {32'hc1cf5cf6, 32'h417e4bb8} /* (3, 1, 14) {real, imag} */,
  {32'h423e5143, 32'hc1389732} /* (3, 1, 13) {real, imag} */,
  {32'hc24ca7c8, 32'h4236d2aa} /* (3, 1, 12) {real, imag} */,
  {32'h416275d2, 32'h41ca126e} /* (3, 1, 11) {real, imag} */,
  {32'h429e5cff, 32'h41d4dd10} /* (3, 1, 10) {real, imag} */,
  {32'h4200fe80, 32'h42d32d16} /* (3, 1, 9) {real, imag} */,
  {32'hc29d4c87, 32'h43118d27} /* (3, 1, 8) {real, imag} */,
  {32'h41ac97fc, 32'hc289026a} /* (3, 1, 7) {real, imag} */,
  {32'h41cae78c, 32'hc2a5c8b8} /* (3, 1, 6) {real, imag} */,
  {32'h43019672, 32'h429fca6f} /* (3, 1, 5) {real, imag} */,
  {32'h42ec2c6b, 32'h438620c7} /* (3, 1, 4) {real, imag} */,
  {32'h429dfe6a, 32'h4205c217} /* (3, 1, 3) {real, imag} */,
  {32'hc3b2aa4d, 32'h43fd2d6b} /* (3, 1, 2) {real, imag} */,
  {32'hc41281ab, 32'hc4a143f0} /* (3, 1, 1) {real, imag} */,
  {32'h41089ec4, 32'h00000000} /* (3, 1, 0) {real, imag} */,
  {32'hc4124592, 32'h44561210} /* (3, 0, 31) {real, imag} */,
  {32'hc3047fcc, 32'hc3bd8ba0} /* (3, 0, 30) {real, imag} */,
  {32'h42866d08, 32'hc205acd8} /* (3, 0, 29) {real, imag} */,
  {32'h4272ce60, 32'hc352e882} /* (3, 0, 28) {real, imag} */,
  {32'h432c58cc, 32'h42503e36} /* (3, 0, 27) {real, imag} */,
  {32'h4220aa6e, 32'h41f47164} /* (3, 0, 26) {real, imag} */,
  {32'h424bb656, 32'h3fc5f450} /* (3, 0, 25) {real, imag} */,
  {32'hc185ba4a, 32'hbf9b1bc0} /* (3, 0, 24) {real, imag} */,
  {32'hc29f20c7, 32'hc1ad5c84} /* (3, 0, 23) {real, imag} */,
  {32'hbfc81440, 32'hc10232f2} /* (3, 0, 22) {real, imag} */,
  {32'hc1aba97e, 32'h41c3ecf9} /* (3, 0, 21) {real, imag} */,
  {32'hc1d5cfb5, 32'h42004ff0} /* (3, 0, 20) {real, imag} */,
  {32'hc1b1ac5c, 32'h4051a3c8} /* (3, 0, 19) {real, imag} */,
  {32'h407b15a0, 32'hc29bfc57} /* (3, 0, 18) {real, imag} */,
  {32'h424b082e, 32'hc1a168cb} /* (3, 0, 17) {real, imag} */,
  {32'hc1188870, 32'h00000000} /* (3, 0, 16) {real, imag} */,
  {32'h424b082e, 32'h41a168cb} /* (3, 0, 15) {real, imag} */,
  {32'h407b15a0, 32'h429bfc57} /* (3, 0, 14) {real, imag} */,
  {32'hc1b1ac5c, 32'hc051a3c8} /* (3, 0, 13) {real, imag} */,
  {32'hc1d5cfb5, 32'hc2004ff0} /* (3, 0, 12) {real, imag} */,
  {32'hc1aba97e, 32'hc1c3ecf9} /* (3, 0, 11) {real, imag} */,
  {32'hbfc81440, 32'h410232f2} /* (3, 0, 10) {real, imag} */,
  {32'hc29f20c7, 32'h41ad5c84} /* (3, 0, 9) {real, imag} */,
  {32'hc185ba4a, 32'h3f9b1bc0} /* (3, 0, 8) {real, imag} */,
  {32'h424bb656, 32'hbfc5f450} /* (3, 0, 7) {real, imag} */,
  {32'h4220aa6e, 32'hc1f47164} /* (3, 0, 6) {real, imag} */,
  {32'h432c58cc, 32'hc2503e36} /* (3, 0, 5) {real, imag} */,
  {32'h4272ce60, 32'h4352e882} /* (3, 0, 4) {real, imag} */,
  {32'h42866d08, 32'h4205acd8} /* (3, 0, 3) {real, imag} */,
  {32'hc3047fcc, 32'h43bd8ba0} /* (3, 0, 2) {real, imag} */,
  {32'hc4124592, 32'hc4561210} /* (3, 0, 1) {real, imag} */,
  {32'h434dfa9a, 32'h00000000} /* (3, 0, 0) {real, imag} */,
  {32'hc48b5903, 32'h43c995f0} /* (2, 31, 31) {real, imag} */,
  {32'h43e34841, 32'hc39d9d6e} /* (2, 31, 30) {real, imag} */,
  {32'h42728d0d, 32'h4239d3b0} /* (2, 31, 29) {real, imag} */,
  {32'hc28538c4, 32'hc2d1403e} /* (2, 31, 28) {real, imag} */,
  {32'h42c98b1c, 32'hc29f64b4} /* (2, 31, 27) {real, imag} */,
  {32'hc210e51c, 32'hc2ed4b70} /* (2, 31, 26) {real, imag} */,
  {32'h41e9744a, 32'h3fc3ace0} /* (2, 31, 25) {real, imag} */,
  {32'h42aa4a55, 32'hc2743a42} /* (2, 31, 24) {real, imag} */,
  {32'h424f9148, 32'h41fef4de} /* (2, 31, 23) {real, imag} */,
  {32'h42550dfa, 32'h420bcfa1} /* (2, 31, 22) {real, imag} */,
  {32'hc17bd9d4, 32'hc2e783e9} /* (2, 31, 21) {real, imag} */,
  {32'h410b74a8, 32'hc0d7cda0} /* (2, 31, 20) {real, imag} */,
  {32'h42552d4f, 32'h42031178} /* (2, 31, 19) {real, imag} */,
  {32'hc1e895b5, 32'hc2067566} /* (2, 31, 18) {real, imag} */,
  {32'h423426be, 32'h414850c8} /* (2, 31, 17) {real, imag} */,
  {32'h4264088f, 32'h00000000} /* (2, 31, 16) {real, imag} */,
  {32'h423426be, 32'hc14850c8} /* (2, 31, 15) {real, imag} */,
  {32'hc1e895b5, 32'h42067566} /* (2, 31, 14) {real, imag} */,
  {32'h42552d4f, 32'hc2031178} /* (2, 31, 13) {real, imag} */,
  {32'h410b74a8, 32'h40d7cda0} /* (2, 31, 12) {real, imag} */,
  {32'hc17bd9d4, 32'h42e783e9} /* (2, 31, 11) {real, imag} */,
  {32'h42550dfa, 32'hc20bcfa1} /* (2, 31, 10) {real, imag} */,
  {32'h424f9148, 32'hc1fef4de} /* (2, 31, 9) {real, imag} */,
  {32'h42aa4a55, 32'h42743a42} /* (2, 31, 8) {real, imag} */,
  {32'h41e9744a, 32'hbfc3ace0} /* (2, 31, 7) {real, imag} */,
  {32'hc210e51c, 32'h42ed4b70} /* (2, 31, 6) {real, imag} */,
  {32'h42c98b1c, 32'h429f64b4} /* (2, 31, 5) {real, imag} */,
  {32'hc28538c4, 32'h42d1403e} /* (2, 31, 4) {real, imag} */,
  {32'h42728d0d, 32'hc239d3b0} /* (2, 31, 3) {real, imag} */,
  {32'h43e34841, 32'h439d9d6e} /* (2, 31, 2) {real, imag} */,
  {32'hc48b5903, 32'hc3c995f0} /* (2, 31, 1) {real, imag} */,
  {32'hc3d50de2, 32'h00000000} /* (2, 31, 0) {real, imag} */,
  {32'hc4ba18fc, 32'h436fc7d8} /* (2, 30, 31) {real, imag} */,
  {32'h44408630, 32'hc354ef78} /* (2, 30, 30) {real, imag} */,
  {32'h42c09fd8, 32'hc1d81e3e} /* (2, 30, 29) {real, imag} */,
  {32'hc28e0f71, 32'hc24b3d9c} /* (2, 30, 28) {real, imag} */,
  {32'h436dcb20, 32'hc2be23c7} /* (2, 30, 27) {real, imag} */,
  {32'hc223b794, 32'hc2b72c3c} /* (2, 30, 26) {real, imag} */,
  {32'hc06aaef8, 32'h426fb155} /* (2, 30, 25) {real, imag} */,
  {32'h431a9a38, 32'hc2b02cd4} /* (2, 30, 24) {real, imag} */,
  {32'hc1978379, 32'h415624d3} /* (2, 30, 23) {real, imag} */,
  {32'h42817ada, 32'h42d3133c} /* (2, 30, 22) {real, imag} */,
  {32'h4322901a, 32'hc24e5121} /* (2, 30, 21) {real, imag} */,
  {32'h42b67872, 32'h428a0b86} /* (2, 30, 20) {real, imag} */,
  {32'hbfb4f6e0, 32'h41289e56} /* (2, 30, 19) {real, imag} */,
  {32'hc2b51a30, 32'h4262a1ae} /* (2, 30, 18) {real, imag} */,
  {32'hc28a5c14, 32'h40aff3d4} /* (2, 30, 17) {real, imag} */,
  {32'hc30ec0fc, 32'h00000000} /* (2, 30, 16) {real, imag} */,
  {32'hc28a5c14, 32'hc0aff3d4} /* (2, 30, 15) {real, imag} */,
  {32'hc2b51a30, 32'hc262a1ae} /* (2, 30, 14) {real, imag} */,
  {32'hbfb4f6e0, 32'hc1289e56} /* (2, 30, 13) {real, imag} */,
  {32'h42b67872, 32'hc28a0b86} /* (2, 30, 12) {real, imag} */,
  {32'h4322901a, 32'h424e5121} /* (2, 30, 11) {real, imag} */,
  {32'h42817ada, 32'hc2d3133c} /* (2, 30, 10) {real, imag} */,
  {32'hc1978379, 32'hc15624d3} /* (2, 30, 9) {real, imag} */,
  {32'h431a9a38, 32'h42b02cd4} /* (2, 30, 8) {real, imag} */,
  {32'hc06aaef8, 32'hc26fb155} /* (2, 30, 7) {real, imag} */,
  {32'hc223b794, 32'h42b72c3c} /* (2, 30, 6) {real, imag} */,
  {32'h436dcb20, 32'h42be23c7} /* (2, 30, 5) {real, imag} */,
  {32'hc28e0f71, 32'h424b3d9c} /* (2, 30, 4) {real, imag} */,
  {32'h42c09fd8, 32'h41d81e3e} /* (2, 30, 3) {real, imag} */,
  {32'h44408630, 32'h4354ef78} /* (2, 30, 2) {real, imag} */,
  {32'hc4ba18fc, 32'hc36fc7d8} /* (2, 30, 1) {real, imag} */,
  {32'hc400a990, 32'h00000000} /* (2, 30, 0) {real, imag} */,
  {32'hc4d64dc6, 32'h437b2d58} /* (2, 29, 31) {real, imag} */,
  {32'h4475c000, 32'hc0f21ec0} /* (2, 29, 30) {real, imag} */,
  {32'h42f5f60e, 32'hc3718a87} /* (2, 29, 29) {real, imag} */,
  {32'hc2d1846a, 32'h41c5d9f4} /* (2, 29, 28) {real, imag} */,
  {32'h4393a75b, 32'hc2d71922} /* (2, 29, 27) {real, imag} */,
  {32'hc16c67e0, 32'h4150abe4} /* (2, 29, 26) {real, imag} */,
  {32'h4214e1d8, 32'h41d2013a} /* (2, 29, 25) {real, imag} */,
  {32'h4307c660, 32'hc2a8209e} /* (2, 29, 24) {real, imag} */,
  {32'hc1e9359c, 32'h42b9f0eb} /* (2, 29, 23) {real, imag} */,
  {32'h421e03e0, 32'h419a60b3} /* (2, 29, 22) {real, imag} */,
  {32'hc1f13add, 32'hc230a678} /* (2, 29, 21) {real, imag} */,
  {32'h4014d7a0, 32'h41f698c0} /* (2, 29, 20) {real, imag} */,
  {32'hc1c693ad, 32'h430853ce} /* (2, 29, 19) {real, imag} */,
  {32'h42bccd05, 32'h41f437fe} /* (2, 29, 18) {real, imag} */,
  {32'hc20be510, 32'hc12f35bf} /* (2, 29, 17) {real, imag} */,
  {32'hc2cc1c6b, 32'h00000000} /* (2, 29, 16) {real, imag} */,
  {32'hc20be510, 32'h412f35bf} /* (2, 29, 15) {real, imag} */,
  {32'h42bccd05, 32'hc1f437fe} /* (2, 29, 14) {real, imag} */,
  {32'hc1c693ad, 32'hc30853ce} /* (2, 29, 13) {real, imag} */,
  {32'h4014d7a0, 32'hc1f698c0} /* (2, 29, 12) {real, imag} */,
  {32'hc1f13add, 32'h4230a678} /* (2, 29, 11) {real, imag} */,
  {32'h421e03e0, 32'hc19a60b3} /* (2, 29, 10) {real, imag} */,
  {32'hc1e9359c, 32'hc2b9f0eb} /* (2, 29, 9) {real, imag} */,
  {32'h4307c660, 32'h42a8209e} /* (2, 29, 8) {real, imag} */,
  {32'h4214e1d8, 32'hc1d2013a} /* (2, 29, 7) {real, imag} */,
  {32'hc16c67e0, 32'hc150abe4} /* (2, 29, 6) {real, imag} */,
  {32'h4393a75b, 32'h42d71922} /* (2, 29, 5) {real, imag} */,
  {32'hc2d1846a, 32'hc1c5d9f4} /* (2, 29, 4) {real, imag} */,
  {32'h42f5f60e, 32'h43718a87} /* (2, 29, 3) {real, imag} */,
  {32'h4475c000, 32'h40f21ec0} /* (2, 29, 2) {real, imag} */,
  {32'hc4d64dc6, 32'hc37b2d58} /* (2, 29, 1) {real, imag} */,
  {32'hc41325e4, 32'h00000000} /* (2, 29, 0) {real, imag} */,
  {32'hc4ecfb29, 32'h42f6a888} /* (2, 28, 31) {real, imag} */,
  {32'h448d2378, 32'h421d8a2a} /* (2, 28, 30) {real, imag} */,
  {32'h428291f3, 32'hc305f861} /* (2, 28, 29) {real, imag} */,
  {32'hc305b184, 32'h430cb0d8} /* (2, 28, 28) {real, imag} */,
  {32'h43a8f5a4, 32'hc33655b4} /* (2, 28, 27) {real, imag} */,
  {32'h4161e0a6, 32'hc10c04f0} /* (2, 28, 26) {real, imag} */,
  {32'hc29d1894, 32'h433c7d9d} /* (2, 28, 25) {real, imag} */,
  {32'h4296c092, 32'h42291555} /* (2, 28, 24) {real, imag} */,
  {32'hc29f0158, 32'hc28f8a09} /* (2, 28, 23) {real, imag} */,
  {32'hc12f0429, 32'h40cd5e90} /* (2, 28, 22) {real, imag} */,
  {32'h42736f61, 32'hc2303064} /* (2, 28, 21) {real, imag} */,
  {32'h42a4ac29, 32'h41bf34e8} /* (2, 28, 20) {real, imag} */,
  {32'h4120e8e0, 32'h4255339a} /* (2, 28, 19) {real, imag} */,
  {32'h41edee1d, 32'h40e627fe} /* (2, 28, 18) {real, imag} */,
  {32'hc25ad449, 32'hc28b8da4} /* (2, 28, 17) {real, imag} */,
  {32'h42648277, 32'h00000000} /* (2, 28, 16) {real, imag} */,
  {32'hc25ad449, 32'h428b8da4} /* (2, 28, 15) {real, imag} */,
  {32'h41edee1d, 32'hc0e627fe} /* (2, 28, 14) {real, imag} */,
  {32'h4120e8e0, 32'hc255339a} /* (2, 28, 13) {real, imag} */,
  {32'h42a4ac29, 32'hc1bf34e8} /* (2, 28, 12) {real, imag} */,
  {32'h42736f61, 32'h42303064} /* (2, 28, 11) {real, imag} */,
  {32'hc12f0429, 32'hc0cd5e90} /* (2, 28, 10) {real, imag} */,
  {32'hc29f0158, 32'h428f8a09} /* (2, 28, 9) {real, imag} */,
  {32'h4296c092, 32'hc2291555} /* (2, 28, 8) {real, imag} */,
  {32'hc29d1894, 32'hc33c7d9d} /* (2, 28, 7) {real, imag} */,
  {32'h4161e0a6, 32'h410c04f0} /* (2, 28, 6) {real, imag} */,
  {32'h43a8f5a4, 32'h433655b4} /* (2, 28, 5) {real, imag} */,
  {32'hc305b184, 32'hc30cb0d8} /* (2, 28, 4) {real, imag} */,
  {32'h428291f3, 32'h4305f861} /* (2, 28, 3) {real, imag} */,
  {32'h448d2378, 32'hc21d8a2a} /* (2, 28, 2) {real, imag} */,
  {32'hc4ecfb29, 32'hc2f6a888} /* (2, 28, 1) {real, imag} */,
  {32'hc42b9c34, 32'h00000000} /* (2, 28, 0) {real, imag} */,
  {32'hc4f64b7e, 32'h42fa6c90} /* (2, 27, 31) {real, imag} */,
  {32'h44797d96, 32'hc2cd985f} /* (2, 27, 30) {real, imag} */,
  {32'h430425b8, 32'hc32d09e8} /* (2, 27, 29) {real, imag} */,
  {32'hc3345c40, 32'h421a704d} /* (2, 27, 28) {real, imag} */,
  {32'h435f5e1a, 32'hc330c00c} /* (2, 27, 27) {real, imag} */,
  {32'hc1dc4b69, 32'hc1b48a16} /* (2, 27, 26) {real, imag} */,
  {32'h418d30aa, 32'h4214d1ea} /* (2, 27, 25) {real, imag} */,
  {32'h4344bd1e, 32'hc1b298dd} /* (2, 27, 24) {real, imag} */,
  {32'h41f453c8, 32'h422e4d2a} /* (2, 27, 23) {real, imag} */,
  {32'h4293ced9, 32'h41bd261f} /* (2, 27, 22) {real, imag} */,
  {32'h40002820, 32'hc215e6e4} /* (2, 27, 21) {real, imag} */,
  {32'h41648678, 32'h42bcced9} /* (2, 27, 20) {real, imag} */,
  {32'hc2d9f0ff, 32'h4228aba6} /* (2, 27, 19) {real, imag} */,
  {32'hc2c4975f, 32'hc1e52c58} /* (2, 27, 18) {real, imag} */,
  {32'hc0abd578, 32'h40c9fefc} /* (2, 27, 17) {real, imag} */,
  {32'hc2bb3816, 32'h00000000} /* (2, 27, 16) {real, imag} */,
  {32'hc0abd578, 32'hc0c9fefc} /* (2, 27, 15) {real, imag} */,
  {32'hc2c4975f, 32'h41e52c58} /* (2, 27, 14) {real, imag} */,
  {32'hc2d9f0ff, 32'hc228aba6} /* (2, 27, 13) {real, imag} */,
  {32'h41648678, 32'hc2bcced9} /* (2, 27, 12) {real, imag} */,
  {32'h40002820, 32'h4215e6e4} /* (2, 27, 11) {real, imag} */,
  {32'h4293ced9, 32'hc1bd261f} /* (2, 27, 10) {real, imag} */,
  {32'h41f453c8, 32'hc22e4d2a} /* (2, 27, 9) {real, imag} */,
  {32'h4344bd1e, 32'h41b298dd} /* (2, 27, 8) {real, imag} */,
  {32'h418d30aa, 32'hc214d1ea} /* (2, 27, 7) {real, imag} */,
  {32'hc1dc4b69, 32'h41b48a16} /* (2, 27, 6) {real, imag} */,
  {32'h435f5e1a, 32'h4330c00c} /* (2, 27, 5) {real, imag} */,
  {32'hc3345c40, 32'hc21a704d} /* (2, 27, 4) {real, imag} */,
  {32'h430425b8, 32'h432d09e8} /* (2, 27, 3) {real, imag} */,
  {32'h44797d96, 32'h42cd985f} /* (2, 27, 2) {real, imag} */,
  {32'hc4f64b7e, 32'hc2fa6c90} /* (2, 27, 1) {real, imag} */,
  {32'hc41a3520, 32'h00000000} /* (2, 27, 0) {real, imag} */,
  {32'hc4f90fbb, 32'h43592860} /* (2, 26, 31) {real, imag} */,
  {32'h44550220, 32'hc25d00f4} /* (2, 26, 30) {real, imag} */,
  {32'h42f31d94, 32'hc2c24364} /* (2, 26, 29) {real, imag} */,
  {32'hc389fc3c, 32'h42261cf2} /* (2, 26, 28) {real, imag} */,
  {32'h4366c6ec, 32'hc2e7c840} /* (2, 26, 27) {real, imag} */,
  {32'h41fd18ce, 32'hc2c366a9} /* (2, 26, 26) {real, imag} */,
  {32'hc2520d71, 32'hc277a026} /* (2, 26, 25) {real, imag} */,
  {32'h430a2718, 32'h41ceb9a5} /* (2, 26, 24) {real, imag} */,
  {32'hc142eb8a, 32'h420beadd} /* (2, 26, 23) {real, imag} */,
  {32'h4200d20c, 32'h42f8bed8} /* (2, 26, 22) {real, imag} */,
  {32'h42706023, 32'hc26cf621} /* (2, 26, 21) {real, imag} */,
  {32'hbf4dc6c0, 32'hc10b6d10} /* (2, 26, 20) {real, imag} */,
  {32'h42b5a7bd, 32'hc2e5ebec} /* (2, 26, 19) {real, imag} */,
  {32'hc1aa705f, 32'h42103a86} /* (2, 26, 18) {real, imag} */,
  {32'hc26c005f, 32'h3fccc590} /* (2, 26, 17) {real, imag} */,
  {32'h42a87456, 32'h00000000} /* (2, 26, 16) {real, imag} */,
  {32'hc26c005f, 32'hbfccc590} /* (2, 26, 15) {real, imag} */,
  {32'hc1aa705f, 32'hc2103a86} /* (2, 26, 14) {real, imag} */,
  {32'h42b5a7bd, 32'h42e5ebec} /* (2, 26, 13) {real, imag} */,
  {32'hbf4dc6c0, 32'h410b6d10} /* (2, 26, 12) {real, imag} */,
  {32'h42706023, 32'h426cf621} /* (2, 26, 11) {real, imag} */,
  {32'h4200d20c, 32'hc2f8bed8} /* (2, 26, 10) {real, imag} */,
  {32'hc142eb8a, 32'hc20beadd} /* (2, 26, 9) {real, imag} */,
  {32'h430a2718, 32'hc1ceb9a5} /* (2, 26, 8) {real, imag} */,
  {32'hc2520d71, 32'h4277a026} /* (2, 26, 7) {real, imag} */,
  {32'h41fd18ce, 32'h42c366a9} /* (2, 26, 6) {real, imag} */,
  {32'h4366c6ec, 32'h42e7c840} /* (2, 26, 5) {real, imag} */,
  {32'hc389fc3c, 32'hc2261cf2} /* (2, 26, 4) {real, imag} */,
  {32'h42f31d94, 32'h42c24364} /* (2, 26, 3) {real, imag} */,
  {32'h44550220, 32'h425d00f4} /* (2, 26, 2) {real, imag} */,
  {32'hc4f90fbb, 32'hc3592860} /* (2, 26, 1) {real, imag} */,
  {32'hc3e7416e, 32'h00000000} /* (2, 26, 0) {real, imag} */,
  {32'hc5003bbd, 32'h432f920c} /* (2, 25, 31) {real, imag} */,
  {32'h44634fac, 32'hc27a4a7a} /* (2, 25, 30) {real, imag} */,
  {32'h42b65f2c, 32'hc2e28299} /* (2, 25, 29) {real, imag} */,
  {32'hc3a9c8e6, 32'h42ad6016} /* (2, 25, 28) {real, imag} */,
  {32'h42ce57d4, 32'hc2807738} /* (2, 25, 27) {real, imag} */,
  {32'h4237a780, 32'hc2aca2a5} /* (2, 25, 26) {real, imag} */,
  {32'hc1d99f08, 32'h429cb5ce} /* (2, 25, 25) {real, imag} */,
  {32'h41c1e119, 32'hc2d477f2} /* (2, 25, 24) {real, imag} */,
  {32'h42d73bcc, 32'h41655a18} /* (2, 25, 23) {real, imag} */,
  {32'hc289c7d3, 32'h42e7cd40} /* (2, 25, 22) {real, imag} */,
  {32'h42545d51, 32'hc2928e7c} /* (2, 25, 21) {real, imag} */,
  {32'hc28c3086, 32'hc250e904} /* (2, 25, 20) {real, imag} */,
  {32'hc2da92c1, 32'h3ef0c700} /* (2, 25, 19) {real, imag} */,
  {32'hc18d441a, 32'hc1907e7a} /* (2, 25, 18) {real, imag} */,
  {32'hc2588ec4, 32'h416c9c50} /* (2, 25, 17) {real, imag} */,
  {32'hc248845d, 32'h00000000} /* (2, 25, 16) {real, imag} */,
  {32'hc2588ec4, 32'hc16c9c50} /* (2, 25, 15) {real, imag} */,
  {32'hc18d441a, 32'h41907e7a} /* (2, 25, 14) {real, imag} */,
  {32'hc2da92c1, 32'hbef0c700} /* (2, 25, 13) {real, imag} */,
  {32'hc28c3086, 32'h4250e904} /* (2, 25, 12) {real, imag} */,
  {32'h42545d51, 32'h42928e7c} /* (2, 25, 11) {real, imag} */,
  {32'hc289c7d3, 32'hc2e7cd40} /* (2, 25, 10) {real, imag} */,
  {32'h42d73bcc, 32'hc1655a18} /* (2, 25, 9) {real, imag} */,
  {32'h41c1e119, 32'h42d477f2} /* (2, 25, 8) {real, imag} */,
  {32'hc1d99f08, 32'hc29cb5ce} /* (2, 25, 7) {real, imag} */,
  {32'h4237a780, 32'h42aca2a5} /* (2, 25, 6) {real, imag} */,
  {32'h42ce57d4, 32'h42807738} /* (2, 25, 5) {real, imag} */,
  {32'hc3a9c8e6, 32'hc2ad6016} /* (2, 25, 4) {real, imag} */,
  {32'h42b65f2c, 32'h42e28299} /* (2, 25, 3) {real, imag} */,
  {32'h44634fac, 32'h427a4a7a} /* (2, 25, 2) {real, imag} */,
  {32'hc5003bbd, 32'hc32f920c} /* (2, 25, 1) {real, imag} */,
  {32'hc418c7d9, 32'h00000000} /* (2, 25, 0) {real, imag} */,
  {32'hc4f82a5d, 32'h422f9b14} /* (2, 24, 31) {real, imag} */,
  {32'h444fba2c, 32'h42256cd0} /* (2, 24, 30) {real, imag} */,
  {32'h4180a906, 32'hc335876c} /* (2, 24, 29) {real, imag} */,
  {32'hc37c12c2, 32'hc0a6b2e0} /* (2, 24, 28) {real, imag} */,
  {32'h42efa661, 32'hc2ec054e} /* (2, 24, 27) {real, imag} */,
  {32'hc2639d5e, 32'h426f44d5} /* (2, 24, 26) {real, imag} */,
  {32'hc26ccab8, 32'hc197a788} /* (2, 24, 25) {real, imag} */,
  {32'h434343e3, 32'hc245f767} /* (2, 24, 24) {real, imag} */,
  {32'h41e82cbe, 32'h41e84ca1} /* (2, 24, 23) {real, imag} */,
  {32'hc2bfc672, 32'hc1cf30b4} /* (2, 24, 22) {real, imag} */,
  {32'h429dd1d0, 32'hc202281c} /* (2, 24, 21) {real, imag} */,
  {32'h423ba2eb, 32'hc218c0c5} /* (2, 24, 20) {real, imag} */,
  {32'hc255bd40, 32'h4286e9ea} /* (2, 24, 19) {real, imag} */,
  {32'h3f801360, 32'hc2875463} /* (2, 24, 18) {real, imag} */,
  {32'h423ecd66, 32'hc2696c0b} /* (2, 24, 17) {real, imag} */,
  {32'h41f2eb33, 32'h00000000} /* (2, 24, 16) {real, imag} */,
  {32'h423ecd66, 32'h42696c0b} /* (2, 24, 15) {real, imag} */,
  {32'h3f801360, 32'h42875463} /* (2, 24, 14) {real, imag} */,
  {32'hc255bd40, 32'hc286e9ea} /* (2, 24, 13) {real, imag} */,
  {32'h423ba2eb, 32'h4218c0c5} /* (2, 24, 12) {real, imag} */,
  {32'h429dd1d0, 32'h4202281c} /* (2, 24, 11) {real, imag} */,
  {32'hc2bfc672, 32'h41cf30b4} /* (2, 24, 10) {real, imag} */,
  {32'h41e82cbe, 32'hc1e84ca1} /* (2, 24, 9) {real, imag} */,
  {32'h434343e3, 32'h4245f767} /* (2, 24, 8) {real, imag} */,
  {32'hc26ccab8, 32'h4197a788} /* (2, 24, 7) {real, imag} */,
  {32'hc2639d5e, 32'hc26f44d5} /* (2, 24, 6) {real, imag} */,
  {32'h42efa661, 32'h42ec054e} /* (2, 24, 5) {real, imag} */,
  {32'hc37c12c2, 32'h40a6b2e0} /* (2, 24, 4) {real, imag} */,
  {32'h4180a906, 32'h4335876c} /* (2, 24, 3) {real, imag} */,
  {32'h444fba2c, 32'hc2256cd0} /* (2, 24, 2) {real, imag} */,
  {32'hc4f82a5d, 32'hc22f9b14} /* (2, 24, 1) {real, imag} */,
  {32'hc4414f50, 32'h00000000} /* (2, 24, 0) {real, imag} */,
  {32'hc4de55de, 32'h422d4ea4} /* (2, 23, 31) {real, imag} */,
  {32'h4423fb19, 32'h4274597e} /* (2, 23, 30) {real, imag} */,
  {32'hc25bdbd0, 32'hc2d1b60e} /* (2, 23, 29) {real, imag} */,
  {32'hc357c014, 32'h418afe38} /* (2, 23, 28) {real, imag} */,
  {32'h42fe002e, 32'hc36d3ff2} /* (2, 23, 27) {real, imag} */,
  {32'hc1662854, 32'hc0fd5a34} /* (2, 23, 26) {real, imag} */,
  {32'hc1e5ef49, 32'hc2162d58} /* (2, 23, 25) {real, imag} */,
  {32'h42758a50, 32'hc2f138b4} /* (2, 23, 24) {real, imag} */,
  {32'h42376254, 32'hc32020e0} /* (2, 23, 23) {real, imag} */,
  {32'hc21b872f, 32'h4225cdc0} /* (2, 23, 22) {real, imag} */,
  {32'h4257bf8d, 32'hc312e28c} /* (2, 23, 21) {real, imag} */,
  {32'h42725586, 32'h422d13da} /* (2, 23, 20) {real, imag} */,
  {32'h425adbb2, 32'h42254c22} /* (2, 23, 19) {real, imag} */,
  {32'hc183a022, 32'h420be862} /* (2, 23, 18) {real, imag} */,
  {32'h42e85dae, 32'h40587a00} /* (2, 23, 17) {real, imag} */,
  {32'h4260bb50, 32'h00000000} /* (2, 23, 16) {real, imag} */,
  {32'h42e85dae, 32'hc0587a00} /* (2, 23, 15) {real, imag} */,
  {32'hc183a022, 32'hc20be862} /* (2, 23, 14) {real, imag} */,
  {32'h425adbb2, 32'hc2254c22} /* (2, 23, 13) {real, imag} */,
  {32'h42725586, 32'hc22d13da} /* (2, 23, 12) {real, imag} */,
  {32'h4257bf8d, 32'h4312e28c} /* (2, 23, 11) {real, imag} */,
  {32'hc21b872f, 32'hc225cdc0} /* (2, 23, 10) {real, imag} */,
  {32'h42376254, 32'h432020e0} /* (2, 23, 9) {real, imag} */,
  {32'h42758a50, 32'h42f138b4} /* (2, 23, 8) {real, imag} */,
  {32'hc1e5ef49, 32'h42162d58} /* (2, 23, 7) {real, imag} */,
  {32'hc1662854, 32'h40fd5a34} /* (2, 23, 6) {real, imag} */,
  {32'h42fe002e, 32'h436d3ff2} /* (2, 23, 5) {real, imag} */,
  {32'hc357c014, 32'hc18afe38} /* (2, 23, 4) {real, imag} */,
  {32'hc25bdbd0, 32'h42d1b60e} /* (2, 23, 3) {real, imag} */,
  {32'h4423fb19, 32'hc274597e} /* (2, 23, 2) {real, imag} */,
  {32'hc4de55de, 32'hc22d4ea4} /* (2, 23, 1) {real, imag} */,
  {32'hc40cacc7, 32'h00000000} /* (2, 23, 0) {real, imag} */,
  {32'hc4a9d95a, 32'hc126a7d0} /* (2, 22, 31) {real, imag} */,
  {32'h440dae01, 32'hc1ec6178} /* (2, 22, 30) {real, imag} */,
  {32'hc294a4e4, 32'h430f4463} /* (2, 22, 29) {real, imag} */,
  {32'hc3499d8b, 32'hc1e4f424} /* (2, 22, 28) {real, imag} */,
  {32'h43478f3a, 32'hc32881af} /* (2, 22, 27) {real, imag} */,
  {32'hc299fe32, 32'h41b08350} /* (2, 22, 26) {real, imag} */,
  {32'h424c0a8c, 32'h421b7832} /* (2, 22, 25) {real, imag} */,
  {32'hc2618dfc, 32'hc29fd098} /* (2, 22, 24) {real, imag} */,
  {32'hc19cc198, 32'h422fb4ab} /* (2, 22, 23) {real, imag} */,
  {32'h42b613cc, 32'h3f5d8400} /* (2, 22, 22) {real, imag} */,
  {32'hc2b8d642, 32'hc26df531} /* (2, 22, 21) {real, imag} */,
  {32'hc3091f16, 32'h42bfb556} /* (2, 22, 20) {real, imag} */,
  {32'hc285f37a, 32'hc1c5cbbe} /* (2, 22, 19) {real, imag} */,
  {32'h41ebbd55, 32'hc1b53b0e} /* (2, 22, 18) {real, imag} */,
  {32'hc2265c22, 32'h427c463e} /* (2, 22, 17) {real, imag} */,
  {32'h41d01c10, 32'h00000000} /* (2, 22, 16) {real, imag} */,
  {32'hc2265c22, 32'hc27c463e} /* (2, 22, 15) {real, imag} */,
  {32'h41ebbd55, 32'h41b53b0e} /* (2, 22, 14) {real, imag} */,
  {32'hc285f37a, 32'h41c5cbbe} /* (2, 22, 13) {real, imag} */,
  {32'hc3091f16, 32'hc2bfb556} /* (2, 22, 12) {real, imag} */,
  {32'hc2b8d642, 32'h426df531} /* (2, 22, 11) {real, imag} */,
  {32'h42b613cc, 32'hbf5d8400} /* (2, 22, 10) {real, imag} */,
  {32'hc19cc198, 32'hc22fb4ab} /* (2, 22, 9) {real, imag} */,
  {32'hc2618dfc, 32'h429fd098} /* (2, 22, 8) {real, imag} */,
  {32'h424c0a8c, 32'hc21b7832} /* (2, 22, 7) {real, imag} */,
  {32'hc299fe32, 32'hc1b08350} /* (2, 22, 6) {real, imag} */,
  {32'h43478f3a, 32'h432881af} /* (2, 22, 5) {real, imag} */,
  {32'hc3499d8b, 32'h41e4f424} /* (2, 22, 4) {real, imag} */,
  {32'hc294a4e4, 32'hc30f4463} /* (2, 22, 3) {real, imag} */,
  {32'h440dae01, 32'h41ec6178} /* (2, 22, 2) {real, imag} */,
  {32'hc4a9d95a, 32'h4126a7d0} /* (2, 22, 1) {real, imag} */,
  {32'hc3c501ea, 32'h00000000} /* (2, 22, 0) {real, imag} */,
  {32'hc4138ae5, 32'hc2ceda50} /* (2, 21, 31) {real, imag} */,
  {32'h42b914b0, 32'hc200009b} /* (2, 21, 30) {real, imag} */,
  {32'hc2c49330, 32'h41902fe4} /* (2, 21, 29) {real, imag} */,
  {32'hc17dac50, 32'h41d8e346} /* (2, 21, 28) {real, imag} */,
  {32'h41ca807c, 32'hc348f586} /* (2, 21, 27) {real, imag} */,
  {32'h3fd44060, 32'h409168e0} /* (2, 21, 26) {real, imag} */,
  {32'hc1fc0446, 32'h42c4ad44} /* (2, 21, 25) {real, imag} */,
  {32'hc19d4da0, 32'h4187d93e} /* (2, 21, 24) {real, imag} */,
  {32'hc2244bf1, 32'hc1c208c1} /* (2, 21, 23) {real, imag} */,
  {32'h42f9c4f4, 32'h4290ba86} /* (2, 21, 22) {real, imag} */,
  {32'h4102fe90, 32'hc2ecdbd6} /* (2, 21, 21) {real, imag} */,
  {32'h42108346, 32'h41584106} /* (2, 21, 20) {real, imag} */,
  {32'hc2240b6e, 32'h41f8619e} /* (2, 21, 19) {real, imag} */,
  {32'h42326026, 32'hc205bb6d} /* (2, 21, 18) {real, imag} */,
  {32'hc1c1b7ef, 32'h4187e687} /* (2, 21, 17) {real, imag} */,
  {32'h41e5a811, 32'h00000000} /* (2, 21, 16) {real, imag} */,
  {32'hc1c1b7ef, 32'hc187e687} /* (2, 21, 15) {real, imag} */,
  {32'h42326026, 32'h4205bb6d} /* (2, 21, 14) {real, imag} */,
  {32'hc2240b6e, 32'hc1f8619e} /* (2, 21, 13) {real, imag} */,
  {32'h42108346, 32'hc1584106} /* (2, 21, 12) {real, imag} */,
  {32'h4102fe90, 32'h42ecdbd6} /* (2, 21, 11) {real, imag} */,
  {32'h42f9c4f4, 32'hc290ba86} /* (2, 21, 10) {real, imag} */,
  {32'hc2244bf1, 32'h41c208c1} /* (2, 21, 9) {real, imag} */,
  {32'hc19d4da0, 32'hc187d93e} /* (2, 21, 8) {real, imag} */,
  {32'hc1fc0446, 32'hc2c4ad44} /* (2, 21, 7) {real, imag} */,
  {32'h3fd44060, 32'hc09168e0} /* (2, 21, 6) {real, imag} */,
  {32'h41ca807c, 32'h4348f586} /* (2, 21, 5) {real, imag} */,
  {32'hc17dac50, 32'hc1d8e346} /* (2, 21, 4) {real, imag} */,
  {32'hc2c49330, 32'hc1902fe4} /* (2, 21, 3) {real, imag} */,
  {32'h42b914b0, 32'h4200009b} /* (2, 21, 2) {real, imag} */,
  {32'hc4138ae5, 32'h42ceda50} /* (2, 21, 1) {real, imag} */,
  {32'h428ab888, 32'h00000000} /* (2, 21, 0) {real, imag} */,
  {32'h442dec8d, 32'hc3a943e1} /* (2, 20, 31) {real, imag} */,
  {32'hc402f12b, 32'h4297af58} /* (2, 20, 30) {real, imag} */,
  {32'hc34603ba, 32'hc114f602} /* (2, 20, 29) {real, imag} */,
  {32'h4237cb54, 32'hc1dff3c6} /* (2, 20, 28) {real, imag} */,
  {32'hc30b0db2, 32'hc2911e8f} /* (2, 20, 27) {real, imag} */,
  {32'h4050d0a0, 32'h42922b8c} /* (2, 20, 26) {real, imag} */,
  {32'hbf5da420, 32'h42acdefa} /* (2, 20, 25) {real, imag} */,
  {32'h40906bea, 32'h42d9c80e} /* (2, 20, 24) {real, imag} */,
  {32'hc1e5c19d, 32'h40e7b954} /* (2, 20, 23) {real, imag} */,
  {32'h40001118, 32'hc33f1014} /* (2, 20, 22) {real, imag} */,
  {32'hc24f4f2e, 32'h42bb78b6} /* (2, 20, 21) {real, imag} */,
  {32'hc15a5924, 32'h42232210} /* (2, 20, 20) {real, imag} */,
  {32'h4205ad32, 32'h42897ea8} /* (2, 20, 19) {real, imag} */,
  {32'h428046da, 32'hc25a9960} /* (2, 20, 18) {real, imag} */,
  {32'h42176a84, 32'h40afeab2} /* (2, 20, 17) {real, imag} */,
  {32'h409bcda0, 32'h00000000} /* (2, 20, 16) {real, imag} */,
  {32'h42176a84, 32'hc0afeab2} /* (2, 20, 15) {real, imag} */,
  {32'h428046da, 32'h425a9960} /* (2, 20, 14) {real, imag} */,
  {32'h4205ad32, 32'hc2897ea8} /* (2, 20, 13) {real, imag} */,
  {32'hc15a5924, 32'hc2232210} /* (2, 20, 12) {real, imag} */,
  {32'hc24f4f2e, 32'hc2bb78b6} /* (2, 20, 11) {real, imag} */,
  {32'h40001118, 32'h433f1014} /* (2, 20, 10) {real, imag} */,
  {32'hc1e5c19d, 32'hc0e7b954} /* (2, 20, 9) {real, imag} */,
  {32'h40906bea, 32'hc2d9c80e} /* (2, 20, 8) {real, imag} */,
  {32'hbf5da420, 32'hc2acdefa} /* (2, 20, 7) {real, imag} */,
  {32'h4050d0a0, 32'hc2922b8c} /* (2, 20, 6) {real, imag} */,
  {32'hc30b0db2, 32'h42911e8f} /* (2, 20, 5) {real, imag} */,
  {32'h4237cb54, 32'h41dff3c6} /* (2, 20, 4) {real, imag} */,
  {32'hc34603ba, 32'h4114f602} /* (2, 20, 3) {real, imag} */,
  {32'hc402f12b, 32'hc297af58} /* (2, 20, 2) {real, imag} */,
  {32'h442dec8d, 32'h43a943e1} /* (2, 20, 1) {real, imag} */,
  {32'h44466964, 32'h00000000} /* (2, 20, 0) {real, imag} */,
  {32'h44a1774f, 32'hc3be1754} /* (2, 19, 31) {real, imag} */,
  {32'hc448bd10, 32'h4115ab98} /* (2, 19, 30) {real, imag} */,
  {32'hc2c6135e, 32'h43046cb4} /* (2, 19, 29) {real, imag} */,
  {32'h432cf01f, 32'hc28b41b1} /* (2, 19, 28) {real, imag} */,
  {32'hc344f50d, 32'h428a1d5f} /* (2, 19, 27) {real, imag} */,
  {32'hc20e5d02, 32'h423fab80} /* (2, 19, 26) {real, imag} */,
  {32'h418c47a8, 32'h424c9d52} /* (2, 19, 25) {real, imag} */,
  {32'hc09e3400, 32'hc15c6720} /* (2, 19, 24) {real, imag} */,
  {32'hc1de8e8c, 32'hc3006ce9} /* (2, 19, 23) {real, imag} */,
  {32'hc1e89904, 32'hc24e1807} /* (2, 19, 22) {real, imag} */,
  {32'hc31f15bc, 32'h411a74e0} /* (2, 19, 21) {real, imag} */,
  {32'h418e1640, 32'h41f281ad} /* (2, 19, 20) {real, imag} */,
  {32'h412d1986, 32'hc2af036c} /* (2, 19, 19) {real, imag} */,
  {32'hc251beb4, 32'h429ffac8} /* (2, 19, 18) {real, imag} */,
  {32'hc13fefa8, 32'h4198077e} /* (2, 19, 17) {real, imag} */,
  {32'h42462c37, 32'h00000000} /* (2, 19, 16) {real, imag} */,
  {32'hc13fefa8, 32'hc198077e} /* (2, 19, 15) {real, imag} */,
  {32'hc251beb4, 32'hc29ffac8} /* (2, 19, 14) {real, imag} */,
  {32'h412d1986, 32'h42af036c} /* (2, 19, 13) {real, imag} */,
  {32'h418e1640, 32'hc1f281ad} /* (2, 19, 12) {real, imag} */,
  {32'hc31f15bc, 32'hc11a74e0} /* (2, 19, 11) {real, imag} */,
  {32'hc1e89904, 32'h424e1807} /* (2, 19, 10) {real, imag} */,
  {32'hc1de8e8c, 32'h43006ce9} /* (2, 19, 9) {real, imag} */,
  {32'hc09e3400, 32'h415c6720} /* (2, 19, 8) {real, imag} */,
  {32'h418c47a8, 32'hc24c9d52} /* (2, 19, 7) {real, imag} */,
  {32'hc20e5d02, 32'hc23fab80} /* (2, 19, 6) {real, imag} */,
  {32'hc344f50d, 32'hc28a1d5f} /* (2, 19, 5) {real, imag} */,
  {32'h432cf01f, 32'h428b41b1} /* (2, 19, 4) {real, imag} */,
  {32'hc2c6135e, 32'hc3046cb4} /* (2, 19, 3) {real, imag} */,
  {32'hc448bd10, 32'hc115ab98} /* (2, 19, 2) {real, imag} */,
  {32'h44a1774f, 32'h43be1754} /* (2, 19, 1) {real, imag} */,
  {32'h44909813, 32'h00000000} /* (2, 19, 0) {real, imag} */,
  {32'h44c78701, 32'hc3996ed0} /* (2, 18, 31) {real, imag} */,
  {32'hc45ab0ea, 32'hc1a80910} /* (2, 18, 30) {real, imag} */,
  {32'hc327faca, 32'h4281ac5c} /* (2, 18, 29) {real, imag} */,
  {32'h4369408c, 32'hc2a3f7e0} /* (2, 18, 28) {real, imag} */,
  {32'hc30aa292, 32'h433c3ff1} /* (2, 18, 27) {real, imag} */,
  {32'hc2300c28, 32'hc1fb95c3} /* (2, 18, 26) {real, imag} */,
  {32'h3dad5300, 32'hc2337d34} /* (2, 18, 25) {real, imag} */,
  {32'hc27e0d3a, 32'h42b3cc8d} /* (2, 18, 24) {real, imag} */,
  {32'hc060d766, 32'h40e71797} /* (2, 18, 23) {real, imag} */,
  {32'h402df800, 32'h4234a267} /* (2, 18, 22) {real, imag} */,
  {32'hc318a243, 32'h40de4122} /* (2, 18, 21) {real, imag} */,
  {32'hc27ade6e, 32'hc2164d91} /* (2, 18, 20) {real, imag} */,
  {32'h422af93f, 32'hc204d9ac} /* (2, 18, 19) {real, imag} */,
  {32'h42114321, 32'h427d0192} /* (2, 18, 18) {real, imag} */,
  {32'h421734e2, 32'hc1c047ad} /* (2, 18, 17) {real, imag} */,
  {32'hc0249440, 32'h00000000} /* (2, 18, 16) {real, imag} */,
  {32'h421734e2, 32'h41c047ad} /* (2, 18, 15) {real, imag} */,
  {32'h42114321, 32'hc27d0192} /* (2, 18, 14) {real, imag} */,
  {32'h422af93f, 32'h4204d9ac} /* (2, 18, 13) {real, imag} */,
  {32'hc27ade6e, 32'h42164d91} /* (2, 18, 12) {real, imag} */,
  {32'hc318a243, 32'hc0de4122} /* (2, 18, 11) {real, imag} */,
  {32'h402df800, 32'hc234a267} /* (2, 18, 10) {real, imag} */,
  {32'hc060d766, 32'hc0e71797} /* (2, 18, 9) {real, imag} */,
  {32'hc27e0d3a, 32'hc2b3cc8d} /* (2, 18, 8) {real, imag} */,
  {32'h3dad5300, 32'h42337d34} /* (2, 18, 7) {real, imag} */,
  {32'hc2300c28, 32'h41fb95c3} /* (2, 18, 6) {real, imag} */,
  {32'hc30aa292, 32'hc33c3ff1} /* (2, 18, 5) {real, imag} */,
  {32'h4369408c, 32'h42a3f7e0} /* (2, 18, 4) {real, imag} */,
  {32'hc327faca, 32'hc281ac5c} /* (2, 18, 3) {real, imag} */,
  {32'hc45ab0ea, 32'h41a80910} /* (2, 18, 2) {real, imag} */,
  {32'h44c78701, 32'h43996ed0} /* (2, 18, 1) {real, imag} */,
  {32'h448f053e, 32'h00000000} /* (2, 18, 0) {real, imag} */,
  {32'h44d86287, 32'hc36e8093} /* (2, 17, 31) {real, imag} */,
  {32'hc475082a, 32'h42e49f38} /* (2, 17, 30) {real, imag} */,
  {32'h402ae4b0, 32'hc1a247af} /* (2, 17, 29) {real, imag} */,
  {32'h42c255b7, 32'hc3657edd} /* (2, 17, 28) {real, imag} */,
  {32'hc2859522, 32'h4310f6aa} /* (2, 17, 27) {real, imag} */,
  {32'h419b74dc, 32'h3e8895e0} /* (2, 17, 26) {real, imag} */,
  {32'h4146e49e, 32'h42731701} /* (2, 17, 25) {real, imag} */,
  {32'hc28b888e, 32'hc27791ef} /* (2, 17, 24) {real, imag} */,
  {32'hc196f035, 32'h42d0f829} /* (2, 17, 23) {real, imag} */,
  {32'h42b7b442, 32'hc2bc7b87} /* (2, 17, 22) {real, imag} */,
  {32'h42bcefe4, 32'h4299e201} /* (2, 17, 21) {real, imag} */,
  {32'h40d79440, 32'h413f5c98} /* (2, 17, 20) {real, imag} */,
  {32'hbe96c280, 32'h40d51116} /* (2, 17, 19) {real, imag} */,
  {32'h423fb16d, 32'hc2bb9e40} /* (2, 17, 18) {real, imag} */,
  {32'hc2034ac2, 32'hc1ac7a10} /* (2, 17, 17) {real, imag} */,
  {32'h41497d40, 32'h00000000} /* (2, 17, 16) {real, imag} */,
  {32'hc2034ac2, 32'h41ac7a10} /* (2, 17, 15) {real, imag} */,
  {32'h423fb16d, 32'h42bb9e40} /* (2, 17, 14) {real, imag} */,
  {32'hbe96c280, 32'hc0d51116} /* (2, 17, 13) {real, imag} */,
  {32'h40d79440, 32'hc13f5c98} /* (2, 17, 12) {real, imag} */,
  {32'h42bcefe4, 32'hc299e201} /* (2, 17, 11) {real, imag} */,
  {32'h42b7b442, 32'h42bc7b87} /* (2, 17, 10) {real, imag} */,
  {32'hc196f035, 32'hc2d0f829} /* (2, 17, 9) {real, imag} */,
  {32'hc28b888e, 32'h427791ef} /* (2, 17, 8) {real, imag} */,
  {32'h4146e49e, 32'hc2731701} /* (2, 17, 7) {real, imag} */,
  {32'h419b74dc, 32'hbe8895e0} /* (2, 17, 6) {real, imag} */,
  {32'hc2859522, 32'hc310f6aa} /* (2, 17, 5) {real, imag} */,
  {32'h42c255b7, 32'h43657edd} /* (2, 17, 4) {real, imag} */,
  {32'h402ae4b0, 32'h41a247af} /* (2, 17, 3) {real, imag} */,
  {32'hc475082a, 32'hc2e49f38} /* (2, 17, 2) {real, imag} */,
  {32'h44d86287, 32'h436e8093} /* (2, 17, 1) {real, imag} */,
  {32'h448ea7b3, 32'h00000000} /* (2, 17, 0) {real, imag} */,
  {32'h44e14996, 32'hc3587a34} /* (2, 16, 31) {real, imag} */,
  {32'hc461adae, 32'h43240e60} /* (2, 16, 30) {real, imag} */,
  {32'h42b08626, 32'h427bb436} /* (2, 16, 29) {real, imag} */,
  {32'h435b42b1, 32'hc30d230d} /* (2, 16, 28) {real, imag} */,
  {32'hc31a1e2e, 32'h42a7d12f} /* (2, 16, 27) {real, imag} */,
  {32'hc125d8d2, 32'h423b030b} /* (2, 16, 26) {real, imag} */,
  {32'h40d2e618, 32'hc2ec8a38} /* (2, 16, 25) {real, imag} */,
  {32'hc3258804, 32'h4193f2c0} /* (2, 16, 24) {real, imag} */,
  {32'h4111f9ea, 32'hc2bdc523} /* (2, 16, 23) {real, imag} */,
  {32'h423d19c0, 32'hc29def97} /* (2, 16, 22) {real, imag} */,
  {32'h40459c80, 32'hc1d9cf30} /* (2, 16, 21) {real, imag} */,
  {32'h4281a096, 32'hc239cba9} /* (2, 16, 20) {real, imag} */,
  {32'h4193596b, 32'h420f449c} /* (2, 16, 19) {real, imag} */,
  {32'hc1883dd4, 32'h42cb642e} /* (2, 16, 18) {real, imag} */,
  {32'h41860f3e, 32'h400b9370} /* (2, 16, 17) {real, imag} */,
  {32'h4201d1a0, 32'h00000000} /* (2, 16, 16) {real, imag} */,
  {32'h41860f3e, 32'hc00b9370} /* (2, 16, 15) {real, imag} */,
  {32'hc1883dd4, 32'hc2cb642e} /* (2, 16, 14) {real, imag} */,
  {32'h4193596b, 32'hc20f449c} /* (2, 16, 13) {real, imag} */,
  {32'h4281a096, 32'h4239cba9} /* (2, 16, 12) {real, imag} */,
  {32'h40459c80, 32'h41d9cf30} /* (2, 16, 11) {real, imag} */,
  {32'h423d19c0, 32'h429def97} /* (2, 16, 10) {real, imag} */,
  {32'h4111f9ea, 32'h42bdc523} /* (2, 16, 9) {real, imag} */,
  {32'hc3258804, 32'hc193f2c0} /* (2, 16, 8) {real, imag} */,
  {32'h40d2e618, 32'h42ec8a38} /* (2, 16, 7) {real, imag} */,
  {32'hc125d8d2, 32'hc23b030b} /* (2, 16, 6) {real, imag} */,
  {32'hc31a1e2e, 32'hc2a7d12f} /* (2, 16, 5) {real, imag} */,
  {32'h435b42b1, 32'h430d230d} /* (2, 16, 4) {real, imag} */,
  {32'h42b08626, 32'hc27bb436} /* (2, 16, 3) {real, imag} */,
  {32'hc461adae, 32'hc3240e60} /* (2, 16, 2) {real, imag} */,
  {32'h44e14996, 32'h43587a34} /* (2, 16, 1) {real, imag} */,
  {32'h44a2e624, 32'h00000000} /* (2, 16, 0) {real, imag} */,
  {32'h44e1a4cd, 32'hc38458c8} /* (2, 15, 31) {real, imag} */,
  {32'hc44a9112, 32'h430a2c30} /* (2, 15, 30) {real, imag} */,
  {32'h4282965e, 32'hc2126220} /* (2, 15, 29) {real, imag} */,
  {32'h432e0488, 32'hc2deb526} /* (2, 15, 28) {real, imag} */,
  {32'hc32d48c2, 32'h4320cea0} /* (2, 15, 27) {real, imag} */,
  {32'hc2d08703, 32'h40c71d7e} /* (2, 15, 26) {real, imag} */,
  {32'h4093831c, 32'hc28b0f0e} /* (2, 15, 25) {real, imag} */,
  {32'hc144769c, 32'hc209e0c9} /* (2, 15, 24) {real, imag} */,
  {32'h424a5bee, 32'h418374e8} /* (2, 15, 23) {real, imag} */,
  {32'hc22efcac, 32'hc219e48e} /* (2, 15, 22) {real, imag} */,
  {32'hc3097bc2, 32'h4237794c} /* (2, 15, 21) {real, imag} */,
  {32'hc1d05494, 32'hc2aa7308} /* (2, 15, 20) {real, imag} */,
  {32'hc20bbaec, 32'hc17a1027} /* (2, 15, 19) {real, imag} */,
  {32'hc1e50aee, 32'h41f44122} /* (2, 15, 18) {real, imag} */,
  {32'h4033fd20, 32'h422331a8} /* (2, 15, 17) {real, imag} */,
  {32'h423d945a, 32'h00000000} /* (2, 15, 16) {real, imag} */,
  {32'h4033fd20, 32'hc22331a8} /* (2, 15, 15) {real, imag} */,
  {32'hc1e50aee, 32'hc1f44122} /* (2, 15, 14) {real, imag} */,
  {32'hc20bbaec, 32'h417a1027} /* (2, 15, 13) {real, imag} */,
  {32'hc1d05494, 32'h42aa7308} /* (2, 15, 12) {real, imag} */,
  {32'hc3097bc2, 32'hc237794c} /* (2, 15, 11) {real, imag} */,
  {32'hc22efcac, 32'h4219e48e} /* (2, 15, 10) {real, imag} */,
  {32'h424a5bee, 32'hc18374e8} /* (2, 15, 9) {real, imag} */,
  {32'hc144769c, 32'h4209e0c9} /* (2, 15, 8) {real, imag} */,
  {32'h4093831c, 32'h428b0f0e} /* (2, 15, 7) {real, imag} */,
  {32'hc2d08703, 32'hc0c71d7e} /* (2, 15, 6) {real, imag} */,
  {32'hc32d48c2, 32'hc320cea0} /* (2, 15, 5) {real, imag} */,
  {32'h432e0488, 32'h42deb526} /* (2, 15, 4) {real, imag} */,
  {32'h4282965e, 32'h42126220} /* (2, 15, 3) {real, imag} */,
  {32'hc44a9112, 32'hc30a2c30} /* (2, 15, 2) {real, imag} */,
  {32'h44e1a4cd, 32'h438458c8} /* (2, 15, 1) {real, imag} */,
  {32'h44a1d59d, 32'h00000000} /* (2, 15, 0) {real, imag} */,
  {32'h44f2d2b1, 32'hc35e6264} /* (2, 14, 31) {real, imag} */,
  {32'hc4512bce, 32'h42f9f698} /* (2, 14, 30) {real, imag} */,
  {32'h42eb75fd, 32'hc28a9628} /* (2, 14, 29) {real, imag} */,
  {32'h431d2fe8, 32'hc1497b84} /* (2, 14, 28) {real, imag} */,
  {32'hc37986d4, 32'h435d0f53} /* (2, 14, 27) {real, imag} */,
  {32'hc278cf16, 32'h3ff7b2d0} /* (2, 14, 26) {real, imag} */,
  {32'hc2248442, 32'hc2457a22} /* (2, 14, 25) {real, imag} */,
  {32'hc2d9637d, 32'h41a7d9c4} /* (2, 14, 24) {real, imag} */,
  {32'hc198b1b3, 32'h40a3ff5b} /* (2, 14, 23) {real, imag} */,
  {32'hc21b83e7, 32'hc2a8ca14} /* (2, 14, 22) {real, imag} */,
  {32'h41d6e04a, 32'h41b8b9de} /* (2, 14, 21) {real, imag} */,
  {32'hc235e926, 32'hc2ec8aac} /* (2, 14, 20) {real, imag} */,
  {32'h428c85be, 32'h420fc854} /* (2, 14, 19) {real, imag} */,
  {32'hc277e7c3, 32'hbdf7e100} /* (2, 14, 18) {real, imag} */,
  {32'hc19670a7, 32'hc1d961ad} /* (2, 14, 17) {real, imag} */,
  {32'hc20cd594, 32'h00000000} /* (2, 14, 16) {real, imag} */,
  {32'hc19670a7, 32'h41d961ad} /* (2, 14, 15) {real, imag} */,
  {32'hc277e7c3, 32'h3df7e100} /* (2, 14, 14) {real, imag} */,
  {32'h428c85be, 32'hc20fc854} /* (2, 14, 13) {real, imag} */,
  {32'hc235e926, 32'h42ec8aac} /* (2, 14, 12) {real, imag} */,
  {32'h41d6e04a, 32'hc1b8b9de} /* (2, 14, 11) {real, imag} */,
  {32'hc21b83e7, 32'h42a8ca14} /* (2, 14, 10) {real, imag} */,
  {32'hc198b1b3, 32'hc0a3ff5b} /* (2, 14, 9) {real, imag} */,
  {32'hc2d9637d, 32'hc1a7d9c4} /* (2, 14, 8) {real, imag} */,
  {32'hc2248442, 32'h42457a22} /* (2, 14, 7) {real, imag} */,
  {32'hc278cf16, 32'hbff7b2d0} /* (2, 14, 6) {real, imag} */,
  {32'hc37986d4, 32'hc35d0f53} /* (2, 14, 5) {real, imag} */,
  {32'h431d2fe8, 32'h41497b84} /* (2, 14, 4) {real, imag} */,
  {32'h42eb75fd, 32'h428a9628} /* (2, 14, 3) {real, imag} */,
  {32'hc4512bce, 32'hc2f9f698} /* (2, 14, 2) {real, imag} */,
  {32'h44f2d2b1, 32'h435e6264} /* (2, 14, 1) {real, imag} */,
  {32'h44ae4e76, 32'h00000000} /* (2, 14, 0) {real, imag} */,
  {32'h44e99c5f, 32'hc3da7c8a} /* (2, 13, 31) {real, imag} */,
  {32'hc4531050, 32'hc1c0e28c} /* (2, 13, 30) {real, imag} */,
  {32'h4281a766, 32'hc2ceb8db} /* (2, 13, 29) {real, imag} */,
  {32'h42ee80c2, 32'hc316498a} /* (2, 13, 28) {real, imag} */,
  {32'hc36e6127, 32'h423e2a50} /* (2, 13, 27) {real, imag} */,
  {32'hc1812afc, 32'h42df92d8} /* (2, 13, 26) {real, imag} */,
  {32'h4200e178, 32'h42403058} /* (2, 13, 25) {real, imag} */,
  {32'hc2b0e4ae, 32'h42964a28} /* (2, 13, 24) {real, imag} */,
  {32'h411c4c28, 32'h42d2c533} /* (2, 13, 23) {real, imag} */,
  {32'h4292024f, 32'hc24c72e1} /* (2, 13, 22) {real, imag} */,
  {32'h417a79e0, 32'h41b82e2c} /* (2, 13, 21) {real, imag} */,
  {32'hc1da4d64, 32'hc1de1671} /* (2, 13, 20) {real, imag} */,
  {32'h425bd464, 32'hc030b6c0} /* (2, 13, 19) {real, imag} */,
  {32'hc2b7e8c8, 32'h42c69adc} /* (2, 13, 18) {real, imag} */,
  {32'h41cb9f7e, 32'h41b3a178} /* (2, 13, 17) {real, imag} */,
  {32'h42768361, 32'h00000000} /* (2, 13, 16) {real, imag} */,
  {32'h41cb9f7e, 32'hc1b3a178} /* (2, 13, 15) {real, imag} */,
  {32'hc2b7e8c8, 32'hc2c69adc} /* (2, 13, 14) {real, imag} */,
  {32'h425bd464, 32'h4030b6c0} /* (2, 13, 13) {real, imag} */,
  {32'hc1da4d64, 32'h41de1671} /* (2, 13, 12) {real, imag} */,
  {32'h417a79e0, 32'hc1b82e2c} /* (2, 13, 11) {real, imag} */,
  {32'h4292024f, 32'h424c72e1} /* (2, 13, 10) {real, imag} */,
  {32'h411c4c28, 32'hc2d2c533} /* (2, 13, 9) {real, imag} */,
  {32'hc2b0e4ae, 32'hc2964a28} /* (2, 13, 8) {real, imag} */,
  {32'h4200e178, 32'hc2403058} /* (2, 13, 7) {real, imag} */,
  {32'hc1812afc, 32'hc2df92d8} /* (2, 13, 6) {real, imag} */,
  {32'hc36e6127, 32'hc23e2a50} /* (2, 13, 5) {real, imag} */,
  {32'h42ee80c2, 32'h4316498a} /* (2, 13, 4) {real, imag} */,
  {32'h4281a766, 32'h42ceb8db} /* (2, 13, 3) {real, imag} */,
  {32'hc4531050, 32'h41c0e28c} /* (2, 13, 2) {real, imag} */,
  {32'h44e99c5f, 32'h43da7c8a} /* (2, 13, 1) {real, imag} */,
  {32'h44acf92f, 32'h00000000} /* (2, 13, 0) {real, imag} */,
  {32'h44cdae8a, 32'hc3a7eb6d} /* (2, 12, 31) {real, imag} */,
  {32'hc42b54e9, 32'h42b83836} /* (2, 12, 30) {real, imag} */,
  {32'hc0f23490, 32'h425b8602} /* (2, 12, 29) {real, imag} */,
  {32'h431bfa46, 32'hc2b8d382} /* (2, 12, 28) {real, imag} */,
  {32'hc3283882, 32'h42ae4a65} /* (2, 12, 27) {real, imag} */,
  {32'hc3036fe6, 32'h432a967a} /* (2, 12, 26) {real, imag} */,
  {32'h420e86f6, 32'h42853138} /* (2, 12, 25) {real, imag} */,
  {32'h3ff78be8, 32'h427575dc} /* (2, 12, 24) {real, imag} */,
  {32'h3f76b6e0, 32'hc25ba55c} /* (2, 12, 23) {real, imag} */,
  {32'h420ca32a, 32'hc0aa6ad0} /* (2, 12, 22) {real, imag} */,
  {32'hc2a7d089, 32'hc16fc8b0} /* (2, 12, 21) {real, imag} */,
  {32'h425eeca1, 32'hc00595e8} /* (2, 12, 20) {real, imag} */,
  {32'h406eec24, 32'h42a10c64} /* (2, 12, 19) {real, imag} */,
  {32'h42082289, 32'hc1ac26a8} /* (2, 12, 18) {real, imag} */,
  {32'h41b095c4, 32'hc09b1552} /* (2, 12, 17) {real, imag} */,
  {32'hc236878b, 32'h00000000} /* (2, 12, 16) {real, imag} */,
  {32'h41b095c4, 32'h409b1552} /* (2, 12, 15) {real, imag} */,
  {32'h42082289, 32'h41ac26a8} /* (2, 12, 14) {real, imag} */,
  {32'h406eec24, 32'hc2a10c64} /* (2, 12, 13) {real, imag} */,
  {32'h425eeca1, 32'h400595e8} /* (2, 12, 12) {real, imag} */,
  {32'hc2a7d089, 32'h416fc8b0} /* (2, 12, 11) {real, imag} */,
  {32'h420ca32a, 32'h40aa6ad0} /* (2, 12, 10) {real, imag} */,
  {32'h3f76b6e0, 32'h425ba55c} /* (2, 12, 9) {real, imag} */,
  {32'h3ff78be8, 32'hc27575dc} /* (2, 12, 8) {real, imag} */,
  {32'h420e86f6, 32'hc2853138} /* (2, 12, 7) {real, imag} */,
  {32'hc3036fe6, 32'hc32a967a} /* (2, 12, 6) {real, imag} */,
  {32'hc3283882, 32'hc2ae4a65} /* (2, 12, 5) {real, imag} */,
  {32'h431bfa46, 32'h42b8d382} /* (2, 12, 4) {real, imag} */,
  {32'hc0f23490, 32'hc25b8602} /* (2, 12, 3) {real, imag} */,
  {32'hc42b54e9, 32'hc2b83836} /* (2, 12, 2) {real, imag} */,
  {32'h44cdae8a, 32'h43a7eb6d} /* (2, 12, 1) {real, imag} */,
  {32'h44886524, 32'h00000000} /* (2, 12, 0) {real, imag} */,
  {32'h448dec80, 32'hc2add5b8} /* (2, 11, 31) {real, imag} */,
  {32'hc4015805, 32'h431ee94e} /* (2, 11, 30) {real, imag} */,
  {32'hc25317cf, 32'hc33708c4} /* (2, 11, 29) {real, imag} */,
  {32'h4329a35a, 32'hc3019700} /* (2, 11, 28) {real, imag} */,
  {32'hc2d36051, 32'h42af42f4} /* (2, 11, 27) {real, imag} */,
  {32'hc2d48cfc, 32'h407b3a40} /* (2, 11, 26) {real, imag} */,
  {32'h42659f47, 32'hc236665b} /* (2, 11, 25) {real, imag} */,
  {32'h42830c02, 32'h42b76cee} /* (2, 11, 24) {real, imag} */,
  {32'h42b1dd5c, 32'hc1936ceb} /* (2, 11, 23) {real, imag} */,
  {32'h428adb62, 32'hc1afdf81} /* (2, 11, 22) {real, imag} */,
  {32'hbf475040, 32'h42c18fbe} /* (2, 11, 21) {real, imag} */,
  {32'hc29840dd, 32'h427dc546} /* (2, 11, 20) {real, imag} */,
  {32'hc13a8a22, 32'h3eb256c0} /* (2, 11, 19) {real, imag} */,
  {32'hc2025356, 32'h41ef0696} /* (2, 11, 18) {real, imag} */,
  {32'h4128b9a6, 32'hc2319636} /* (2, 11, 17) {real, imag} */,
  {32'hc06a77b8, 32'h00000000} /* (2, 11, 16) {real, imag} */,
  {32'h4128b9a6, 32'h42319636} /* (2, 11, 15) {real, imag} */,
  {32'hc2025356, 32'hc1ef0696} /* (2, 11, 14) {real, imag} */,
  {32'hc13a8a22, 32'hbeb256c0} /* (2, 11, 13) {real, imag} */,
  {32'hc29840dd, 32'hc27dc546} /* (2, 11, 12) {real, imag} */,
  {32'hbf475040, 32'hc2c18fbe} /* (2, 11, 11) {real, imag} */,
  {32'h428adb62, 32'h41afdf81} /* (2, 11, 10) {real, imag} */,
  {32'h42b1dd5c, 32'h41936ceb} /* (2, 11, 9) {real, imag} */,
  {32'h42830c02, 32'hc2b76cee} /* (2, 11, 8) {real, imag} */,
  {32'h42659f47, 32'h4236665b} /* (2, 11, 7) {real, imag} */,
  {32'hc2d48cfc, 32'hc07b3a40} /* (2, 11, 6) {real, imag} */,
  {32'hc2d36051, 32'hc2af42f4} /* (2, 11, 5) {real, imag} */,
  {32'h4329a35a, 32'h43019700} /* (2, 11, 4) {real, imag} */,
  {32'hc25317cf, 32'h433708c4} /* (2, 11, 3) {real, imag} */,
  {32'hc4015805, 32'hc31ee94e} /* (2, 11, 2) {real, imag} */,
  {32'h448dec80, 32'h42add5b8} /* (2, 11, 1) {real, imag} */,
  {32'h44168693, 32'h00000000} /* (2, 11, 0) {real, imag} */,
  {32'hc395e368, 32'h415f29b0} /* (2, 10, 31) {real, imag} */,
  {32'h4118a5c0, 32'hc2ff7c46} /* (2, 10, 30) {real, imag} */,
  {32'hc270ca44, 32'hc353a7bd} /* (2, 10, 29) {real, imag} */,
  {32'hc2c8b18a, 32'hc318d050} /* (2, 10, 28) {real, imag} */,
  {32'hc2805a2f, 32'hc2ee5a47} /* (2, 10, 27) {real, imag} */,
  {32'h40e279a8, 32'hc14d2174} /* (2, 10, 26) {real, imag} */,
  {32'h42016bae, 32'hc04d8400} /* (2, 10, 25) {real, imag} */,
  {32'h4127c400, 32'hc1cfae62} /* (2, 10, 24) {real, imag} */,
  {32'hbdf52880, 32'hc307a7f4} /* (2, 10, 23) {real, imag} */,
  {32'hc27f6d34, 32'hc01695e0} /* (2, 10, 22) {real, imag} */,
  {32'h42196003, 32'h40b62618} /* (2, 10, 21) {real, imag} */,
  {32'h4068e380, 32'hc0a70800} /* (2, 10, 20) {real, imag} */,
  {32'h42d20cea, 32'hc2814a7c} /* (2, 10, 19) {real, imag} */,
  {32'h422ccaca, 32'hc2d5d1f0} /* (2, 10, 18) {real, imag} */,
  {32'h423bc89e, 32'h40050888} /* (2, 10, 17) {real, imag} */,
  {32'hc2680d88, 32'h00000000} /* (2, 10, 16) {real, imag} */,
  {32'h423bc89e, 32'hc0050888} /* (2, 10, 15) {real, imag} */,
  {32'h422ccaca, 32'h42d5d1f0} /* (2, 10, 14) {real, imag} */,
  {32'h42d20cea, 32'h42814a7c} /* (2, 10, 13) {real, imag} */,
  {32'h4068e380, 32'h40a70800} /* (2, 10, 12) {real, imag} */,
  {32'h42196003, 32'hc0b62618} /* (2, 10, 11) {real, imag} */,
  {32'hc27f6d34, 32'h401695e0} /* (2, 10, 10) {real, imag} */,
  {32'hbdf52880, 32'h4307a7f4} /* (2, 10, 9) {real, imag} */,
  {32'h4127c400, 32'h41cfae62} /* (2, 10, 8) {real, imag} */,
  {32'h42016bae, 32'h404d8400} /* (2, 10, 7) {real, imag} */,
  {32'h40e279a8, 32'h414d2174} /* (2, 10, 6) {real, imag} */,
  {32'hc2805a2f, 32'h42ee5a47} /* (2, 10, 5) {real, imag} */,
  {32'hc2c8b18a, 32'h4318d050} /* (2, 10, 4) {real, imag} */,
  {32'hc270ca44, 32'h4353a7bd} /* (2, 10, 3) {real, imag} */,
  {32'h4118a5c0, 32'h42ff7c46} /* (2, 10, 2) {real, imag} */,
  {32'hc395e368, 32'hc15f29b0} /* (2, 10, 1) {real, imag} */,
  {32'hc34ff884, 32'h00000000} /* (2, 10, 0) {real, imag} */,
  {32'hc482dc4e, 32'h4358bc01} /* (2, 9, 31) {real, imag} */,
  {32'h43b98166, 32'hc384c700} /* (2, 9, 30) {real, imag} */,
  {32'h41d64db4, 32'hc345f5dd} /* (2, 9, 29) {real, imag} */,
  {32'hc2b5d0f1, 32'hc261e420} /* (2, 9, 28) {real, imag} */,
  {32'h42df47ea, 32'hc1e0d7c0} /* (2, 9, 27) {real, imag} */,
  {32'h417b74ec, 32'h4257740e} /* (2, 9, 26) {real, imag} */,
  {32'h420c0d7c, 32'h431e9eb6} /* (2, 9, 25) {real, imag} */,
  {32'h430eaa2f, 32'hc29f5462} /* (2, 9, 24) {real, imag} */,
  {32'hc229bc8a, 32'h42c61285} /* (2, 9, 23) {real, imag} */,
  {32'h420dde69, 32'h424a39e8} /* (2, 9, 22) {real, imag} */,
  {32'h4233ad69, 32'h421c7ea7} /* (2, 9, 21) {real, imag} */,
  {32'h40d4b780, 32'hc1958e1f} /* (2, 9, 20) {real, imag} */,
  {32'h4136e948, 32'h413a30e6} /* (2, 9, 19) {real, imag} */,
  {32'h414abb2b, 32'hc24bc524} /* (2, 9, 18) {real, imag} */,
  {32'h426e468c, 32'h4109a49e} /* (2, 9, 17) {real, imag} */,
  {32'hc2ea8262, 32'h00000000} /* (2, 9, 16) {real, imag} */,
  {32'h426e468c, 32'hc109a49e} /* (2, 9, 15) {real, imag} */,
  {32'h414abb2b, 32'h424bc524} /* (2, 9, 14) {real, imag} */,
  {32'h4136e948, 32'hc13a30e6} /* (2, 9, 13) {real, imag} */,
  {32'h40d4b780, 32'h41958e1f} /* (2, 9, 12) {real, imag} */,
  {32'h4233ad69, 32'hc21c7ea7} /* (2, 9, 11) {real, imag} */,
  {32'h420dde69, 32'hc24a39e8} /* (2, 9, 10) {real, imag} */,
  {32'hc229bc8a, 32'hc2c61285} /* (2, 9, 9) {real, imag} */,
  {32'h430eaa2f, 32'h429f5462} /* (2, 9, 8) {real, imag} */,
  {32'h420c0d7c, 32'hc31e9eb6} /* (2, 9, 7) {real, imag} */,
  {32'h417b74ec, 32'hc257740e} /* (2, 9, 6) {real, imag} */,
  {32'h42df47ea, 32'h41e0d7c0} /* (2, 9, 5) {real, imag} */,
  {32'hc2b5d0f1, 32'h4261e420} /* (2, 9, 4) {real, imag} */,
  {32'h41d64db4, 32'h4345f5dd} /* (2, 9, 3) {real, imag} */,
  {32'h43b98166, 32'h4384c700} /* (2, 9, 2) {real, imag} */,
  {32'hc482dc4e, 32'hc358bc01} /* (2, 9, 1) {real, imag} */,
  {32'hc4475199, 32'h00000000} /* (2, 9, 0) {real, imag} */,
  {32'hc4ad4633, 32'h4339539d} /* (2, 8, 31) {real, imag} */,
  {32'h443322b0, 32'hc28393f8} /* (2, 8, 30) {real, imag} */,
  {32'hc2446779, 32'hc2951b40} /* (2, 8, 29) {real, imag} */,
  {32'hc2c800dc, 32'h427eba14} /* (2, 8, 28) {real, imag} */,
  {32'h43592968, 32'hc2839472} /* (2, 8, 27) {real, imag} */,
  {32'h429b1451, 32'h42e7552c} /* (2, 8, 26) {real, imag} */,
  {32'hc0c25794, 32'h433620a5} /* (2, 8, 25) {real, imag} */,
  {32'h42bf205e, 32'hc1a48a1e} /* (2, 8, 24) {real, imag} */,
  {32'h425bf477, 32'h429b6259} /* (2, 8, 23) {real, imag} */,
  {32'h42164847, 32'h41fbae84} /* (2, 8, 22) {real, imag} */,
  {32'hc25beb67, 32'hc2402cbc} /* (2, 8, 21) {real, imag} */,
  {32'h42c2e672, 32'hc17bbccb} /* (2, 8, 20) {real, imag} */,
  {32'hc1fd875f, 32'hc2b608ac} /* (2, 8, 19) {real, imag} */,
  {32'h4033da60, 32'h40c6d334} /* (2, 8, 18) {real, imag} */,
  {32'hc216ca7e, 32'hc24d9621} /* (2, 8, 17) {real, imag} */,
  {32'h418b86df, 32'h00000000} /* (2, 8, 16) {real, imag} */,
  {32'hc216ca7e, 32'h424d9621} /* (2, 8, 15) {real, imag} */,
  {32'h4033da60, 32'hc0c6d334} /* (2, 8, 14) {real, imag} */,
  {32'hc1fd875f, 32'h42b608ac} /* (2, 8, 13) {real, imag} */,
  {32'h42c2e672, 32'h417bbccb} /* (2, 8, 12) {real, imag} */,
  {32'hc25beb67, 32'h42402cbc} /* (2, 8, 11) {real, imag} */,
  {32'h42164847, 32'hc1fbae84} /* (2, 8, 10) {real, imag} */,
  {32'h425bf477, 32'hc29b6259} /* (2, 8, 9) {real, imag} */,
  {32'h42bf205e, 32'h41a48a1e} /* (2, 8, 8) {real, imag} */,
  {32'hc0c25794, 32'hc33620a5} /* (2, 8, 7) {real, imag} */,
  {32'h429b1451, 32'hc2e7552c} /* (2, 8, 6) {real, imag} */,
  {32'h43592968, 32'h42839472} /* (2, 8, 5) {real, imag} */,
  {32'hc2c800dc, 32'hc27eba14} /* (2, 8, 4) {real, imag} */,
  {32'hc2446779, 32'h42951b40} /* (2, 8, 3) {real, imag} */,
  {32'h443322b0, 32'h428393f8} /* (2, 8, 2) {real, imag} */,
  {32'hc4ad4633, 32'hc339539d} /* (2, 8, 1) {real, imag} */,
  {32'hc48991fc, 32'h00000000} /* (2, 8, 0) {real, imag} */,
  {32'hc4c9b112, 32'h43c83912} /* (2, 7, 31) {real, imag} */,
  {32'h444ee35c, 32'hc2406f5a} /* (2, 7, 30) {real, imag} */,
  {32'h42957f00, 32'hc2e54d1f} /* (2, 7, 29) {real, imag} */,
  {32'hc2aef829, 32'hc3201cd4} /* (2, 7, 28) {real, imag} */,
  {32'h43132b18, 32'h422608c8} /* (2, 7, 27) {real, imag} */,
  {32'h42cb5b98, 32'hc2b65e67} /* (2, 7, 26) {real, imag} */,
  {32'hc242a644, 32'hc24ca314} /* (2, 7, 25) {real, imag} */,
  {32'h424e2c10, 32'hc2d78940} /* (2, 7, 24) {real, imag} */,
  {32'hc278e180, 32'hc1a93724} /* (2, 7, 23) {real, imag} */,
  {32'hc2c20f31, 32'h412ed9e0} /* (2, 7, 22) {real, imag} */,
  {32'h4106eb24, 32'hc326eeec} /* (2, 7, 21) {real, imag} */,
  {32'hc305613b, 32'hc18a9be3} /* (2, 7, 20) {real, imag} */,
  {32'h43078fc0, 32'h42df9077} /* (2, 7, 19) {real, imag} */,
  {32'h4200b031, 32'hc28a5118} /* (2, 7, 18) {real, imag} */,
  {32'h41b44004, 32'hc195d424} /* (2, 7, 17) {real, imag} */,
  {32'h42ca90c0, 32'h00000000} /* (2, 7, 16) {real, imag} */,
  {32'h41b44004, 32'h4195d424} /* (2, 7, 15) {real, imag} */,
  {32'h4200b031, 32'h428a5118} /* (2, 7, 14) {real, imag} */,
  {32'h43078fc0, 32'hc2df9077} /* (2, 7, 13) {real, imag} */,
  {32'hc305613b, 32'h418a9be3} /* (2, 7, 12) {real, imag} */,
  {32'h4106eb24, 32'h4326eeec} /* (2, 7, 11) {real, imag} */,
  {32'hc2c20f31, 32'hc12ed9e0} /* (2, 7, 10) {real, imag} */,
  {32'hc278e180, 32'h41a93724} /* (2, 7, 9) {real, imag} */,
  {32'h424e2c10, 32'h42d78940} /* (2, 7, 8) {real, imag} */,
  {32'hc242a644, 32'h424ca314} /* (2, 7, 7) {real, imag} */,
  {32'h42cb5b98, 32'h42b65e67} /* (2, 7, 6) {real, imag} */,
  {32'h43132b18, 32'hc22608c8} /* (2, 7, 5) {real, imag} */,
  {32'hc2aef829, 32'h43201cd4} /* (2, 7, 4) {real, imag} */,
  {32'h42957f00, 32'h42e54d1f} /* (2, 7, 3) {real, imag} */,
  {32'h444ee35c, 32'h42406f5a} /* (2, 7, 2) {real, imag} */,
  {32'hc4c9b112, 32'hc3c83912} /* (2, 7, 1) {real, imag} */,
  {32'hc4a53e92, 32'h00000000} /* (2, 7, 0) {real, imag} */,
  {32'hc4bde0e9, 32'h4448b732} /* (2, 6, 31) {real, imag} */,
  {32'h441ed100, 32'hc2d9a35a} /* (2, 6, 30) {real, imag} */,
  {32'h438da6dd, 32'h420bc094} /* (2, 6, 29) {real, imag} */,
  {32'hc2eaf458, 32'hc31895da} /* (2, 6, 28) {real, imag} */,
  {32'h4303109c, 32'hc2e7bb76} /* (2, 6, 27) {real, imag} */,
  {32'h42d3cdde, 32'h4144fd18} /* (2, 6, 26) {real, imag} */,
  {32'hc24697cd, 32'hbfa57800} /* (2, 6, 25) {real, imag} */,
  {32'h42c50392, 32'hc21337a0} /* (2, 6, 24) {real, imag} */,
  {32'hbff75964, 32'h42408871} /* (2, 6, 23) {real, imag} */,
  {32'h42b59b90, 32'h40dde648} /* (2, 6, 22) {real, imag} */,
  {32'h41986186, 32'hc2110d7d} /* (2, 6, 21) {real, imag} */,
  {32'hc270362a, 32'h42958b68} /* (2, 6, 20) {real, imag} */,
  {32'hc1d8a489, 32'hc20e5495} /* (2, 6, 19) {real, imag} */,
  {32'h41c7127f, 32'h42021b54} /* (2, 6, 18) {real, imag} */,
  {32'hc29c895a, 32'hc1714992} /* (2, 6, 17) {real, imag} */,
  {32'h423f49b4, 32'h00000000} /* (2, 6, 16) {real, imag} */,
  {32'hc29c895a, 32'h41714992} /* (2, 6, 15) {real, imag} */,
  {32'h41c7127f, 32'hc2021b54} /* (2, 6, 14) {real, imag} */,
  {32'hc1d8a489, 32'h420e5495} /* (2, 6, 13) {real, imag} */,
  {32'hc270362a, 32'hc2958b68} /* (2, 6, 12) {real, imag} */,
  {32'h41986186, 32'h42110d7d} /* (2, 6, 11) {real, imag} */,
  {32'h42b59b90, 32'hc0dde648} /* (2, 6, 10) {real, imag} */,
  {32'hbff75964, 32'hc2408871} /* (2, 6, 9) {real, imag} */,
  {32'h42c50392, 32'h421337a0} /* (2, 6, 8) {real, imag} */,
  {32'hc24697cd, 32'h3fa57800} /* (2, 6, 7) {real, imag} */,
  {32'h42d3cdde, 32'hc144fd18} /* (2, 6, 6) {real, imag} */,
  {32'h4303109c, 32'h42e7bb76} /* (2, 6, 5) {real, imag} */,
  {32'hc2eaf458, 32'h431895da} /* (2, 6, 4) {real, imag} */,
  {32'h438da6dd, 32'hc20bc094} /* (2, 6, 3) {real, imag} */,
  {32'h441ed100, 32'h42d9a35a} /* (2, 6, 2) {real, imag} */,
  {32'hc4bde0e9, 32'hc448b732} /* (2, 6, 1) {real, imag} */,
  {32'hc48b89d4, 32'h00000000} /* (2, 6, 0) {real, imag} */,
  {32'hc4967b12, 32'h4495996f} /* (2, 5, 31) {real, imag} */,
  {32'h430d7946, 32'hc3889242} /* (2, 5, 30) {real, imag} */,
  {32'h43ae0444, 32'hc166e338} /* (2, 5, 29) {real, imag} */,
  {32'hc3336e5c, 32'hc2e7ccb8} /* (2, 5, 28) {real, imag} */,
  {32'h4304c706, 32'hbfc75100} /* (2, 5, 27) {real, imag} */,
  {32'hc165add6, 32'h42fa1aa2} /* (2, 5, 26) {real, imag} */,
  {32'hc2a236b2, 32'h419fa9e5} /* (2, 5, 25) {real, imag} */,
  {32'h41bbea28, 32'h42455210} /* (2, 5, 24) {real, imag} */,
  {32'hc216a4ea, 32'h4290a478} /* (2, 5, 23) {real, imag} */,
  {32'hc23f53c2, 32'hc22c6360} /* (2, 5, 22) {real, imag} */,
  {32'h42bc3cf3, 32'hbe5baa00} /* (2, 5, 21) {real, imag} */,
  {32'hbf077fc0, 32'hc1f89724} /* (2, 5, 20) {real, imag} */,
  {32'h420cb5da, 32'h4169d941} /* (2, 5, 19) {real, imag} */,
  {32'hc28e31fb, 32'h4270f648} /* (2, 5, 18) {real, imag} */,
  {32'h42af75aa, 32'h4214f5a2} /* (2, 5, 17) {real, imag} */,
  {32'hc2317fcf, 32'h00000000} /* (2, 5, 16) {real, imag} */,
  {32'h42af75aa, 32'hc214f5a2} /* (2, 5, 15) {real, imag} */,
  {32'hc28e31fb, 32'hc270f648} /* (2, 5, 14) {real, imag} */,
  {32'h420cb5da, 32'hc169d941} /* (2, 5, 13) {real, imag} */,
  {32'hbf077fc0, 32'h41f89724} /* (2, 5, 12) {real, imag} */,
  {32'h42bc3cf3, 32'h3e5baa00} /* (2, 5, 11) {real, imag} */,
  {32'hc23f53c2, 32'h422c6360} /* (2, 5, 10) {real, imag} */,
  {32'hc216a4ea, 32'hc290a478} /* (2, 5, 9) {real, imag} */,
  {32'h41bbea28, 32'hc2455210} /* (2, 5, 8) {real, imag} */,
  {32'hc2a236b2, 32'hc19fa9e5} /* (2, 5, 7) {real, imag} */,
  {32'hc165add6, 32'hc2fa1aa2} /* (2, 5, 6) {real, imag} */,
  {32'h4304c706, 32'h3fc75100} /* (2, 5, 5) {real, imag} */,
  {32'hc3336e5c, 32'h42e7ccb8} /* (2, 5, 4) {real, imag} */,
  {32'h43ae0444, 32'h4166e338} /* (2, 5, 3) {real, imag} */,
  {32'h430d7946, 32'h43889242} /* (2, 5, 2) {real, imag} */,
  {32'hc4967b12, 32'hc495996f} /* (2, 5, 1) {real, imag} */,
  {32'hc48444f0, 32'h00000000} /* (2, 5, 0) {real, imag} */,
  {32'hc47d6f5e, 32'h44de33f6} /* (2, 4, 31) {real, imag} */,
  {32'hc38d8048, 32'hc392136b} /* (2, 4, 30) {real, imag} */,
  {32'h4366ec8c, 32'hc0ae3ba0} /* (2, 4, 29) {real, imag} */,
  {32'hc1f193e8, 32'hc30f416a} /* (2, 4, 28) {real, imag} */,
  {32'h4288ff70, 32'h42998269} /* (2, 4, 27) {real, imag} */,
  {32'h40ecaa7c, 32'h42c2e23d} /* (2, 4, 26) {real, imag} */,
  {32'h4328ab32, 32'h42db92be} /* (2, 4, 25) {real, imag} */,
  {32'hc1270918, 32'hc2b46aea} /* (2, 4, 24) {real, imag} */,
  {32'h42c7cecc, 32'hc0acfdc0} /* (2, 4, 23) {real, imag} */,
  {32'h40ef9b36, 32'hc30a073e} /* (2, 4, 22) {real, imag} */,
  {32'hc0a1d4d8, 32'hc1a66b48} /* (2, 4, 21) {real, imag} */,
  {32'hc2a5846f, 32'hc20d6961} /* (2, 4, 20) {real, imag} */,
  {32'h42951d84, 32'hc1063f3c} /* (2, 4, 19) {real, imag} */,
  {32'hc26b9f2c, 32'h42104d89} /* (2, 4, 18) {real, imag} */,
  {32'h42a1af84, 32'hc22e9e62} /* (2, 4, 17) {real, imag} */,
  {32'hc284d047, 32'h00000000} /* (2, 4, 16) {real, imag} */,
  {32'h42a1af84, 32'h422e9e62} /* (2, 4, 15) {real, imag} */,
  {32'hc26b9f2c, 32'hc2104d89} /* (2, 4, 14) {real, imag} */,
  {32'h42951d84, 32'h41063f3c} /* (2, 4, 13) {real, imag} */,
  {32'hc2a5846f, 32'h420d6961} /* (2, 4, 12) {real, imag} */,
  {32'hc0a1d4d8, 32'h41a66b48} /* (2, 4, 11) {real, imag} */,
  {32'h40ef9b36, 32'h430a073e} /* (2, 4, 10) {real, imag} */,
  {32'h42c7cecc, 32'h40acfdc0} /* (2, 4, 9) {real, imag} */,
  {32'hc1270918, 32'h42b46aea} /* (2, 4, 8) {real, imag} */,
  {32'h4328ab32, 32'hc2db92be} /* (2, 4, 7) {real, imag} */,
  {32'h40ecaa7c, 32'hc2c2e23d} /* (2, 4, 6) {real, imag} */,
  {32'h4288ff70, 32'hc2998269} /* (2, 4, 5) {real, imag} */,
  {32'hc1f193e8, 32'h430f416a} /* (2, 4, 4) {real, imag} */,
  {32'h4366ec8c, 32'h40ae3ba0} /* (2, 4, 3) {real, imag} */,
  {32'hc38d8048, 32'h4392136b} /* (2, 4, 2) {real, imag} */,
  {32'hc47d6f5e, 32'hc4de33f6} /* (2, 4, 1) {real, imag} */,
  {32'hc48cc5ce, 32'h00000000} /* (2, 4, 0) {real, imag} */,
  {32'hc4636f08, 32'h44d837eb} /* (2, 3, 31) {real, imag} */,
  {32'hc3d108c1, 32'hc3f695c7} /* (2, 3, 30) {real, imag} */,
  {32'h4382edaa, 32'h41d4eac8} /* (2, 3, 29) {real, imag} */,
  {32'h418b6622, 32'hc33b67b8} /* (2, 3, 28) {real, imag} */,
  {32'h4330cd5e, 32'h428b2652} /* (2, 3, 27) {real, imag} */,
  {32'h422ecfda, 32'h42cf0082} /* (2, 3, 26) {real, imag} */,
  {32'h42826ba0, 32'h429035cc} /* (2, 3, 25) {real, imag} */,
  {32'hc20d996a, 32'hc245736c} /* (2, 3, 24) {real, imag} */,
  {32'h43456ca4, 32'hc2329082} /* (2, 3, 23) {real, imag} */,
  {32'hc1797aa0, 32'hc1fc59f1} /* (2, 3, 22) {real, imag} */,
  {32'h426960da, 32'hc0f32fd0} /* (2, 3, 21) {real, imag} */,
  {32'hc202bda0, 32'hc22f9a90} /* (2, 3, 20) {real, imag} */,
  {32'hc26dec4c, 32'h4144c840} /* (2, 3, 19) {real, imag} */,
  {32'hc0c7e1d0, 32'hc29f0d7a} /* (2, 3, 18) {real, imag} */,
  {32'hc0503150, 32'hc1934032} /* (2, 3, 17) {real, imag} */,
  {32'h426abc02, 32'h00000000} /* (2, 3, 16) {real, imag} */,
  {32'hc0503150, 32'h41934032} /* (2, 3, 15) {real, imag} */,
  {32'hc0c7e1d0, 32'h429f0d7a} /* (2, 3, 14) {real, imag} */,
  {32'hc26dec4c, 32'hc144c840} /* (2, 3, 13) {real, imag} */,
  {32'hc202bda0, 32'h422f9a90} /* (2, 3, 12) {real, imag} */,
  {32'h426960da, 32'h40f32fd0} /* (2, 3, 11) {real, imag} */,
  {32'hc1797aa0, 32'h41fc59f1} /* (2, 3, 10) {real, imag} */,
  {32'h43456ca4, 32'h42329082} /* (2, 3, 9) {real, imag} */,
  {32'hc20d996a, 32'h4245736c} /* (2, 3, 8) {real, imag} */,
  {32'h42826ba0, 32'hc29035cc} /* (2, 3, 7) {real, imag} */,
  {32'h422ecfda, 32'hc2cf0082} /* (2, 3, 6) {real, imag} */,
  {32'h4330cd5e, 32'hc28b2652} /* (2, 3, 5) {real, imag} */,
  {32'h418b6622, 32'h433b67b8} /* (2, 3, 4) {real, imag} */,
  {32'h4382edaa, 32'hc1d4eac8} /* (2, 3, 3) {real, imag} */,
  {32'hc3d108c1, 32'h43f695c7} /* (2, 3, 2) {real, imag} */,
  {32'hc4636f08, 32'hc4d837eb} /* (2, 3, 1) {real, imag} */,
  {32'hc4701ed4, 32'h00000000} /* (2, 3, 0) {real, imag} */,
  {32'hc45ea864, 32'h44cedacb} /* (2, 2, 31) {real, imag} */,
  {32'hc3e1d8c7, 32'hc44dd26a} /* (2, 2, 30) {real, imag} */,
  {32'h435e7844, 32'h42920072} /* (2, 2, 29) {real, imag} */,
  {32'h433f1150, 32'hc3a26c70} /* (2, 2, 28) {real, imag} */,
  {32'h42a7fe43, 32'h4279c092} /* (2, 2, 27) {real, imag} */,
  {32'h4246656c, 32'h42533ba4} /* (2, 2, 26) {real, imag} */,
  {32'h4266b8c6, 32'hc08eb698} /* (2, 2, 25) {real, imag} */,
  {32'hc2814da1, 32'hc2f3a16e} /* (2, 2, 24) {real, imag} */,
  {32'hc1a2fff3, 32'h414bf4fd} /* (2, 2, 23) {real, imag} */,
  {32'hc19289bf, 32'hc2849128} /* (2, 2, 22) {real, imag} */,
  {32'h417d6360, 32'hc18d3c0e} /* (2, 2, 21) {real, imag} */,
  {32'h4196ddf2, 32'hc1f3ecbb} /* (2, 2, 20) {real, imag} */,
  {32'hc28fa238, 32'hc219fc5a} /* (2, 2, 19) {real, imag} */,
  {32'h42583145, 32'hc2f017a1} /* (2, 2, 18) {real, imag} */,
  {32'h42def736, 32'h42459416} /* (2, 2, 17) {real, imag} */,
  {32'h41e77754, 32'h00000000} /* (2, 2, 16) {real, imag} */,
  {32'h42def736, 32'hc2459416} /* (2, 2, 15) {real, imag} */,
  {32'h42583145, 32'h42f017a1} /* (2, 2, 14) {real, imag} */,
  {32'hc28fa238, 32'h4219fc5a} /* (2, 2, 13) {real, imag} */,
  {32'h4196ddf2, 32'h41f3ecbb} /* (2, 2, 12) {real, imag} */,
  {32'h417d6360, 32'h418d3c0e} /* (2, 2, 11) {real, imag} */,
  {32'hc19289bf, 32'h42849128} /* (2, 2, 10) {real, imag} */,
  {32'hc1a2fff3, 32'hc14bf4fd} /* (2, 2, 9) {real, imag} */,
  {32'hc2814da1, 32'h42f3a16e} /* (2, 2, 8) {real, imag} */,
  {32'h4266b8c6, 32'h408eb698} /* (2, 2, 7) {real, imag} */,
  {32'h4246656c, 32'hc2533ba4} /* (2, 2, 6) {real, imag} */,
  {32'h42a7fe43, 32'hc279c092} /* (2, 2, 5) {real, imag} */,
  {32'h433f1150, 32'h43a26c70} /* (2, 2, 4) {real, imag} */,
  {32'h435e7844, 32'hc2920072} /* (2, 2, 3) {real, imag} */,
  {32'hc3e1d8c7, 32'h444dd26a} /* (2, 2, 2) {real, imag} */,
  {32'hc45ea864, 32'hc4cedacb} /* (2, 2, 1) {real, imag} */,
  {32'hc465f67e, 32'h00000000} /* (2, 2, 0) {real, imag} */,
  {32'hc46c95e2, 32'h44b469fc} /* (2, 1, 31) {real, imag} */,
  {32'hc3b017a3, 32'hc42c29d0} /* (2, 1, 30) {real, imag} */,
  {32'h42ffe39e, 32'hbfe6d810} /* (2, 1, 29) {real, imag} */,
  {32'h4274f81c, 32'hc3985e8c} /* (2, 1, 28) {real, imag} */,
  {32'h4289e2be, 32'h42ba21c8} /* (2, 1, 27) {real, imag} */,
  {32'h41cceed7, 32'h4296314e} /* (2, 1, 26) {real, imag} */,
  {32'hc279db1b, 32'h42be54a8} /* (2, 1, 25) {real, imag} */,
  {32'hc27a6246, 32'h404bd660} /* (2, 1, 24) {real, imag} */,
  {32'hc2a7bb42, 32'hc30450ae} /* (2, 1, 23) {real, imag} */,
  {32'h41b718c5, 32'hc3032ea4} /* (2, 1, 22) {real, imag} */,
  {32'h430558db, 32'hc1569338} /* (2, 1, 21) {real, imag} */,
  {32'h422be5c8, 32'h4213b4d6} /* (2, 1, 20) {real, imag} */,
  {32'h40dd7180, 32'hc184a6bd} /* (2, 1, 19) {real, imag} */,
  {32'hc10a90a6, 32'hbf9b12d0} /* (2, 1, 18) {real, imag} */,
  {32'h41fa81a0, 32'hc222dd12} /* (2, 1, 17) {real, imag} */,
  {32'hc2892994, 32'h00000000} /* (2, 1, 16) {real, imag} */,
  {32'h41fa81a0, 32'h4222dd12} /* (2, 1, 15) {real, imag} */,
  {32'hc10a90a6, 32'h3f9b12d0} /* (2, 1, 14) {real, imag} */,
  {32'h40dd7180, 32'h4184a6bd} /* (2, 1, 13) {real, imag} */,
  {32'h422be5c8, 32'hc213b4d6} /* (2, 1, 12) {real, imag} */,
  {32'h430558db, 32'h41569338} /* (2, 1, 11) {real, imag} */,
  {32'h41b718c5, 32'h43032ea4} /* (2, 1, 10) {real, imag} */,
  {32'hc2a7bb42, 32'h430450ae} /* (2, 1, 9) {real, imag} */,
  {32'hc27a6246, 32'hc04bd660} /* (2, 1, 8) {real, imag} */,
  {32'hc279db1b, 32'hc2be54a8} /* (2, 1, 7) {real, imag} */,
  {32'h41cceed7, 32'hc296314e} /* (2, 1, 6) {real, imag} */,
  {32'h4289e2be, 32'hc2ba21c8} /* (2, 1, 5) {real, imag} */,
  {32'h4274f81c, 32'h43985e8c} /* (2, 1, 4) {real, imag} */,
  {32'h42ffe39e, 32'h3fe6d810} /* (2, 1, 3) {real, imag} */,
  {32'hc3b017a3, 32'h442c29d0} /* (2, 1, 2) {real, imag} */,
  {32'hc46c95e2, 32'hc4b469fc} /* (2, 1, 1) {real, imag} */,
  {32'hc3dd49b2, 32'h00000000} /* (2, 1, 0) {real, imag} */,
  {32'hc45a1c5c, 32'h4472038b} /* (2, 0, 31) {real, imag} */,
  {32'hc2b71410, 32'hc3e25ce0} /* (2, 0, 30) {real, imag} */,
  {32'h41b118e2, 32'hc293e7c7} /* (2, 0, 29) {real, imag} */,
  {32'hc1fdd1c8, 32'hc33a9b03} /* (2, 0, 28) {real, imag} */,
  {32'h4326e388, 32'h41c92c64} /* (2, 0, 27) {real, imag} */,
  {32'h428939a1, 32'h41ae8e92} /* (2, 0, 26) {real, imag} */,
  {32'hc2f9432a, 32'h42751f2d} /* (2, 0, 25) {real, imag} */,
  {32'hc2950453, 32'h421fd9ae} /* (2, 0, 24) {real, imag} */,
  {32'hc1ecb9c5, 32'hc2e869fd} /* (2, 0, 23) {real, imag} */,
  {32'h42c0a5a0, 32'hc2d814ad} /* (2, 0, 22) {real, imag} */,
  {32'h42464faa, 32'h42ade000} /* (2, 0, 21) {real, imag} */,
  {32'h41ef2a66, 32'h422e2ebd} /* (2, 0, 20) {real, imag} */,
  {32'hc2090fb6, 32'hbfa55dd0} /* (2, 0, 19) {real, imag} */,
  {32'hc284a8c1, 32'h40ab6200} /* (2, 0, 18) {real, imag} */,
  {32'hc1340cbb, 32'hc2317a3c} /* (2, 0, 17) {real, imag} */,
  {32'hc0ef11cc, 32'h00000000} /* (2, 0, 16) {real, imag} */,
  {32'hc1340cbb, 32'h42317a3c} /* (2, 0, 15) {real, imag} */,
  {32'hc284a8c1, 32'hc0ab6200} /* (2, 0, 14) {real, imag} */,
  {32'hc2090fb6, 32'h3fa55dd0} /* (2, 0, 13) {real, imag} */,
  {32'h41ef2a66, 32'hc22e2ebd} /* (2, 0, 12) {real, imag} */,
  {32'h42464faa, 32'hc2ade000} /* (2, 0, 11) {real, imag} */,
  {32'h42c0a5a0, 32'h42d814ad} /* (2, 0, 10) {real, imag} */,
  {32'hc1ecb9c5, 32'h42e869fd} /* (2, 0, 9) {real, imag} */,
  {32'hc2950453, 32'hc21fd9ae} /* (2, 0, 8) {real, imag} */,
  {32'hc2f9432a, 32'hc2751f2d} /* (2, 0, 7) {real, imag} */,
  {32'h428939a1, 32'hc1ae8e92} /* (2, 0, 6) {real, imag} */,
  {32'h4326e388, 32'hc1c92c64} /* (2, 0, 5) {real, imag} */,
  {32'hc1fdd1c8, 32'h433a9b03} /* (2, 0, 4) {real, imag} */,
  {32'h41b118e2, 32'h4293e7c7} /* (2, 0, 3) {real, imag} */,
  {32'hc2b71410, 32'h43e25ce0} /* (2, 0, 2) {real, imag} */,
  {32'hc45a1c5c, 32'hc472038b} /* (2, 0, 1) {real, imag} */,
  {32'hc3a3cf8f, 32'h00000000} /* (2, 0, 0) {real, imag} */,
  {32'hc468585e, 32'h43e20071} /* (1, 31, 31) {real, imag} */,
  {32'h43a47fec, 32'hc362088f} /* (1, 31, 30) {real, imag} */,
  {32'h42809d40, 32'h420475b4} /* (1, 31, 29) {real, imag} */,
  {32'h3fef6d30, 32'h41daa6f0} /* (1, 31, 28) {real, imag} */,
  {32'h4336690d, 32'hc1e211fc} /* (1, 31, 27) {real, imag} */,
  {32'hc22b61bc, 32'hc294faf0} /* (1, 31, 26) {real, imag} */,
  {32'hc1af03a8, 32'h41c2b31e} /* (1, 31, 25) {real, imag} */,
  {32'hc217d5b5, 32'hc2c3610a} /* (1, 31, 24) {real, imag} */,
  {32'h418ac1bc, 32'h423a61c4} /* (1, 31, 23) {real, imag} */,
  {32'h4246d4fa, 32'hc1b6db9a} /* (1, 31, 22) {real, imag} */,
  {32'h42a540f6, 32'hc1f2893c} /* (1, 31, 21) {real, imag} */,
  {32'h421e530a, 32'h419a655f} /* (1, 31, 20) {real, imag} */,
  {32'hc20cbab5, 32'h41cbd0f0} /* (1, 31, 19) {real, imag} */,
  {32'h41a3a20e, 32'hc2509d42} /* (1, 31, 18) {real, imag} */,
  {32'hc2083fa9, 32'hc1c6743c} /* (1, 31, 17) {real, imag} */,
  {32'hbff24f00, 32'h00000000} /* (1, 31, 16) {real, imag} */,
  {32'hc2083fa9, 32'h41c6743c} /* (1, 31, 15) {real, imag} */,
  {32'h41a3a20e, 32'h42509d42} /* (1, 31, 14) {real, imag} */,
  {32'hc20cbab5, 32'hc1cbd0f0} /* (1, 31, 13) {real, imag} */,
  {32'h421e530a, 32'hc19a655f} /* (1, 31, 12) {real, imag} */,
  {32'h42a540f6, 32'h41f2893c} /* (1, 31, 11) {real, imag} */,
  {32'h4246d4fa, 32'h41b6db9a} /* (1, 31, 10) {real, imag} */,
  {32'h418ac1bc, 32'hc23a61c4} /* (1, 31, 9) {real, imag} */,
  {32'hc217d5b5, 32'h42c3610a} /* (1, 31, 8) {real, imag} */,
  {32'hc1af03a8, 32'hc1c2b31e} /* (1, 31, 7) {real, imag} */,
  {32'hc22b61bc, 32'h4294faf0} /* (1, 31, 6) {real, imag} */,
  {32'h4336690d, 32'h41e211fc} /* (1, 31, 5) {real, imag} */,
  {32'h3fef6d30, 32'hc1daa6f0} /* (1, 31, 4) {real, imag} */,
  {32'h42809d40, 32'hc20475b4} /* (1, 31, 3) {real, imag} */,
  {32'h43a47fec, 32'h4362088f} /* (1, 31, 2) {real, imag} */,
  {32'hc468585e, 32'hc3e20071} /* (1, 31, 1) {real, imag} */,
  {32'hc4028506, 32'h00000000} /* (1, 31, 0) {real, imag} */,
  {32'hc493059a, 32'h434b15b0} /* (1, 30, 31) {real, imag} */,
  {32'h4416f75b, 32'hc3551c14} /* (1, 30, 30) {real, imag} */,
  {32'h42dd1033, 32'hc0395d20} /* (1, 30, 29) {real, imag} */,
  {32'h42576eca, 32'h42780570} /* (1, 30, 28) {real, imag} */,
  {32'h43020744, 32'hc302f2ad} /* (1, 30, 27) {real, imag} */,
  {32'h41faee26, 32'hc2fc2341} /* (1, 30, 26) {real, imag} */,
  {32'hc3053feb, 32'h42a555b8} /* (1, 30, 25) {real, imag} */,
  {32'h41e2668c, 32'hc24bd587} /* (1, 30, 24) {real, imag} */,
  {32'hc2a260db, 32'h429de8b1} /* (1, 30, 23) {real, imag} */,
  {32'hc28550d2, 32'h4315b2b8} /* (1, 30, 22) {real, imag} */,
  {32'h40d0a060, 32'hc1acb2ae} /* (1, 30, 21) {real, imag} */,
  {32'h4155d47c, 32'hc1e6d732} /* (1, 30, 20) {real, imag} */,
  {32'h406378e8, 32'h4206797a} /* (1, 30, 19) {real, imag} */,
  {32'hc0e24ce8, 32'hc296b4cb} /* (1, 30, 18) {real, imag} */,
  {32'hc297c4a2, 32'h413449ac} /* (1, 30, 17) {real, imag} */,
  {32'h41c59562, 32'h00000000} /* (1, 30, 16) {real, imag} */,
  {32'hc297c4a2, 32'hc13449ac} /* (1, 30, 15) {real, imag} */,
  {32'hc0e24ce8, 32'h4296b4cb} /* (1, 30, 14) {real, imag} */,
  {32'h406378e8, 32'hc206797a} /* (1, 30, 13) {real, imag} */,
  {32'h4155d47c, 32'h41e6d732} /* (1, 30, 12) {real, imag} */,
  {32'h40d0a060, 32'h41acb2ae} /* (1, 30, 11) {real, imag} */,
  {32'hc28550d2, 32'hc315b2b8} /* (1, 30, 10) {real, imag} */,
  {32'hc2a260db, 32'hc29de8b1} /* (1, 30, 9) {real, imag} */,
  {32'h41e2668c, 32'h424bd587} /* (1, 30, 8) {real, imag} */,
  {32'hc3053feb, 32'hc2a555b8} /* (1, 30, 7) {real, imag} */,
  {32'h41faee26, 32'h42fc2341} /* (1, 30, 6) {real, imag} */,
  {32'h43020744, 32'h4302f2ad} /* (1, 30, 5) {real, imag} */,
  {32'h42576eca, 32'hc2780570} /* (1, 30, 4) {real, imag} */,
  {32'h42dd1033, 32'h40395d20} /* (1, 30, 3) {real, imag} */,
  {32'h4416f75b, 32'h43551c14} /* (1, 30, 2) {real, imag} */,
  {32'hc493059a, 32'hc34b15b0} /* (1, 30, 1) {real, imag} */,
  {32'hc423405f, 32'h00000000} /* (1, 30, 0) {real, imag} */,
  {32'hc4b50e2b, 32'h41d0f5c0} /* (1, 29, 31) {real, imag} */,
  {32'h443f7aa2, 32'hc362fb75} /* (1, 29, 30) {real, imag} */,
  {32'h4213721e, 32'hc24538d7} /* (1, 29, 29) {real, imag} */,
  {32'h40aa29d0, 32'h4283b664} /* (1, 29, 28) {real, imag} */,
  {32'h4398464e, 32'hc19b2a80} /* (1, 29, 27) {real, imag} */,
  {32'h4183d7ee, 32'h41366bfa} /* (1, 29, 26) {real, imag} */,
  {32'hc2f582ae, 32'h42ac1a8a} /* (1, 29, 25) {real, imag} */,
  {32'h41d2dc94, 32'hc27eb8bb} /* (1, 29, 24) {real, imag} */,
  {32'hc15d2f18, 32'hc2c029de} /* (1, 29, 23) {real, imag} */,
  {32'hc28d7e25, 32'h424d537e} /* (1, 29, 22) {real, imag} */,
  {32'h423dd078, 32'hc18391d0} /* (1, 29, 21) {real, imag} */,
  {32'h41afd642, 32'h42243957} /* (1, 29, 20) {real, imag} */,
  {32'h40a9be20, 32'h408ccc36} /* (1, 29, 19) {real, imag} */,
  {32'h4199b69e, 32'h4172eea8} /* (1, 29, 18) {real, imag} */,
  {32'hc094a55a, 32'h4191cad6} /* (1, 29, 17) {real, imag} */,
  {32'hc1042fcc, 32'h00000000} /* (1, 29, 16) {real, imag} */,
  {32'hc094a55a, 32'hc191cad6} /* (1, 29, 15) {real, imag} */,
  {32'h4199b69e, 32'hc172eea8} /* (1, 29, 14) {real, imag} */,
  {32'h40a9be20, 32'hc08ccc36} /* (1, 29, 13) {real, imag} */,
  {32'h41afd642, 32'hc2243957} /* (1, 29, 12) {real, imag} */,
  {32'h423dd078, 32'h418391d0} /* (1, 29, 11) {real, imag} */,
  {32'hc28d7e25, 32'hc24d537e} /* (1, 29, 10) {real, imag} */,
  {32'hc15d2f18, 32'h42c029de} /* (1, 29, 9) {real, imag} */,
  {32'h41d2dc94, 32'h427eb8bb} /* (1, 29, 8) {real, imag} */,
  {32'hc2f582ae, 32'hc2ac1a8a} /* (1, 29, 7) {real, imag} */,
  {32'h4183d7ee, 32'hc1366bfa} /* (1, 29, 6) {real, imag} */,
  {32'h4398464e, 32'h419b2a80} /* (1, 29, 5) {real, imag} */,
  {32'h40aa29d0, 32'hc283b664} /* (1, 29, 4) {real, imag} */,
  {32'h4213721e, 32'h424538d7} /* (1, 29, 3) {real, imag} */,
  {32'h443f7aa2, 32'h4362fb75} /* (1, 29, 2) {real, imag} */,
  {32'hc4b50e2b, 32'hc1d0f5c0} /* (1, 29, 1) {real, imag} */,
  {32'hc449ea6b, 32'h00000000} /* (1, 29, 0) {real, imag} */,
  {32'hc4c40ace, 32'h43102880} /* (1, 28, 31) {real, imag} */,
  {32'h443be20a, 32'hc211c0b8} /* (1, 28, 30) {real, imag} */,
  {32'h41fb73d0, 32'hc244409c} /* (1, 28, 29) {real, imag} */,
  {32'hc3362b3b, 32'h4316165d} /* (1, 28, 28) {real, imag} */,
  {32'h436754ad, 32'hc2782426} /* (1, 28, 27) {real, imag} */,
  {32'hc1e9af26, 32'h422443bb} /* (1, 28, 26) {real, imag} */,
  {32'h409a8b30, 32'h427ead96} /* (1, 28, 25) {real, imag} */,
  {32'h42f2bc74, 32'hc2be18ac} /* (1, 28, 24) {real, imag} */,
  {32'hc2bc4a2e, 32'hc1cc6208} /* (1, 28, 23) {real, imag} */,
  {32'hc23c033a, 32'hc2b99ea0} /* (1, 28, 22) {real, imag} */,
  {32'hc1b23e6e, 32'hc282b69d} /* (1, 28, 21) {real, imag} */,
  {32'hc137cefa, 32'h429a552a} /* (1, 28, 20) {real, imag} */,
  {32'hc1dee6a0, 32'h41ad4061} /* (1, 28, 19) {real, imag} */,
  {32'hc152bee8, 32'hc0ff6864} /* (1, 28, 18) {real, imag} */,
  {32'h417621d4, 32'hc1923df5} /* (1, 28, 17) {real, imag} */,
  {32'h4066f6e8, 32'h00000000} /* (1, 28, 16) {real, imag} */,
  {32'h417621d4, 32'h41923df5} /* (1, 28, 15) {real, imag} */,
  {32'hc152bee8, 32'h40ff6864} /* (1, 28, 14) {real, imag} */,
  {32'hc1dee6a0, 32'hc1ad4061} /* (1, 28, 13) {real, imag} */,
  {32'hc137cefa, 32'hc29a552a} /* (1, 28, 12) {real, imag} */,
  {32'hc1b23e6e, 32'h4282b69d} /* (1, 28, 11) {real, imag} */,
  {32'hc23c033a, 32'h42b99ea0} /* (1, 28, 10) {real, imag} */,
  {32'hc2bc4a2e, 32'h41cc6208} /* (1, 28, 9) {real, imag} */,
  {32'h42f2bc74, 32'h42be18ac} /* (1, 28, 8) {real, imag} */,
  {32'h409a8b30, 32'hc27ead96} /* (1, 28, 7) {real, imag} */,
  {32'hc1e9af26, 32'hc22443bb} /* (1, 28, 6) {real, imag} */,
  {32'h436754ad, 32'h42782426} /* (1, 28, 5) {real, imag} */,
  {32'hc3362b3b, 32'hc316165d} /* (1, 28, 4) {real, imag} */,
  {32'h41fb73d0, 32'h4244409c} /* (1, 28, 3) {real, imag} */,
  {32'h443be20a, 32'h4211c0b8} /* (1, 28, 2) {real, imag} */,
  {32'hc4c40ace, 32'hc3102880} /* (1, 28, 1) {real, imag} */,
  {32'hc4460cd1, 32'h00000000} /* (1, 28, 0) {real, imag} */,
  {32'hc4d559aa, 32'h4301d9cc} /* (1, 27, 31) {real, imag} */,
  {32'h4427b2bb, 32'h4250dbf8} /* (1, 27, 30) {real, imag} */,
  {32'h428c4f58, 32'hc29749c3} /* (1, 27, 29) {real, imag} */,
  {32'hc310a81d, 32'h43473848} /* (1, 27, 28) {real, imag} */,
  {32'h43a83587, 32'hc27966f7} /* (1, 27, 27) {real, imag} */,
  {32'h42be8d07, 32'hc2dd6439} /* (1, 27, 26) {real, imag} */,
  {32'h41f68b3a, 32'hc13414b0} /* (1, 27, 25) {real, imag} */,
  {32'h425b6df1, 32'hc2f0e8e6} /* (1, 27, 24) {real, imag} */,
  {32'hc211f298, 32'hc23d341b} /* (1, 27, 23) {real, imag} */,
  {32'hc118470e, 32'h41593c02} /* (1, 27, 22) {real, imag} */,
  {32'h41c1e870, 32'h420aa1f2} /* (1, 27, 21) {real, imag} */,
  {32'hc1a3e1ba, 32'h428f18ae} /* (1, 27, 20) {real, imag} */,
  {32'hc1e18b80, 32'hc2073ef7} /* (1, 27, 19) {real, imag} */,
  {32'hc288c491, 32'hc22dfd2e} /* (1, 27, 18) {real, imag} */,
  {32'hc139fa6a, 32'h428f25f8} /* (1, 27, 17) {real, imag} */,
  {32'h428b913e, 32'h00000000} /* (1, 27, 16) {real, imag} */,
  {32'hc139fa6a, 32'hc28f25f8} /* (1, 27, 15) {real, imag} */,
  {32'hc288c491, 32'h422dfd2e} /* (1, 27, 14) {real, imag} */,
  {32'hc1e18b80, 32'h42073ef7} /* (1, 27, 13) {real, imag} */,
  {32'hc1a3e1ba, 32'hc28f18ae} /* (1, 27, 12) {real, imag} */,
  {32'h41c1e870, 32'hc20aa1f2} /* (1, 27, 11) {real, imag} */,
  {32'hc118470e, 32'hc1593c02} /* (1, 27, 10) {real, imag} */,
  {32'hc211f298, 32'h423d341b} /* (1, 27, 9) {real, imag} */,
  {32'h425b6df1, 32'h42f0e8e6} /* (1, 27, 8) {real, imag} */,
  {32'h41f68b3a, 32'h413414b0} /* (1, 27, 7) {real, imag} */,
  {32'h42be8d07, 32'h42dd6439} /* (1, 27, 6) {real, imag} */,
  {32'h43a83587, 32'h427966f7} /* (1, 27, 5) {real, imag} */,
  {32'hc310a81d, 32'hc3473848} /* (1, 27, 4) {real, imag} */,
  {32'h428c4f58, 32'h429749c3} /* (1, 27, 3) {real, imag} */,
  {32'h4427b2bb, 32'hc250dbf8} /* (1, 27, 2) {real, imag} */,
  {32'hc4d559aa, 32'hc301d9cc} /* (1, 27, 1) {real, imag} */,
  {32'hc411db1a, 32'h00000000} /* (1, 27, 0) {real, imag} */,
  {32'hc4ce6c52, 32'h42ce283a} /* (1, 26, 31) {real, imag} */,
  {32'h4409fd6b, 32'hc170d040} /* (1, 26, 30) {real, imag} */,
  {32'hc24d3202, 32'hc2d30f30} /* (1, 26, 29) {real, imag} */,
  {32'hc305353a, 32'h42a3a4f2} /* (1, 26, 28) {real, imag} */,
  {32'h43624dba, 32'hc30822f9} /* (1, 26, 27) {real, imag} */,
  {32'h430e3c5a, 32'h41f8b26c} /* (1, 26, 26) {real, imag} */,
  {32'hc21066e9, 32'h411e29b0} /* (1, 26, 25) {real, imag} */,
  {32'h42924d57, 32'hc2fb220a} /* (1, 26, 24) {real, imag} */,
  {32'h427b89c4, 32'hc2905d69} /* (1, 26, 23) {real, imag} */,
  {32'hc0eee088, 32'h4266f5b9} /* (1, 26, 22) {real, imag} */,
  {32'hc293261c, 32'hc24ceb08} /* (1, 26, 21) {real, imag} */,
  {32'h41a92f24, 32'hc0914bf8} /* (1, 26, 20) {real, imag} */,
  {32'hc09778c0, 32'hc12d8b14} /* (1, 26, 19) {real, imag} */,
  {32'h40a403b0, 32'h425b3d28} /* (1, 26, 18) {real, imag} */,
  {32'hc17597ae, 32'hc104660c} /* (1, 26, 17) {real, imag} */,
  {32'hc23b56fa, 32'h00000000} /* (1, 26, 16) {real, imag} */,
  {32'hc17597ae, 32'h4104660c} /* (1, 26, 15) {real, imag} */,
  {32'h40a403b0, 32'hc25b3d28} /* (1, 26, 14) {real, imag} */,
  {32'hc09778c0, 32'h412d8b14} /* (1, 26, 13) {real, imag} */,
  {32'h41a92f24, 32'h40914bf8} /* (1, 26, 12) {real, imag} */,
  {32'hc293261c, 32'h424ceb08} /* (1, 26, 11) {real, imag} */,
  {32'hc0eee088, 32'hc266f5b9} /* (1, 26, 10) {real, imag} */,
  {32'h427b89c4, 32'h42905d69} /* (1, 26, 9) {real, imag} */,
  {32'h42924d57, 32'h42fb220a} /* (1, 26, 8) {real, imag} */,
  {32'hc21066e9, 32'hc11e29b0} /* (1, 26, 7) {real, imag} */,
  {32'h430e3c5a, 32'hc1f8b26c} /* (1, 26, 6) {real, imag} */,
  {32'h43624dba, 32'h430822f9} /* (1, 26, 5) {real, imag} */,
  {32'hc305353a, 32'hc2a3a4f2} /* (1, 26, 4) {real, imag} */,
  {32'hc24d3202, 32'h42d30f30} /* (1, 26, 3) {real, imag} */,
  {32'h4409fd6b, 32'h4170d040} /* (1, 26, 2) {real, imag} */,
  {32'hc4ce6c52, 32'hc2ce283a} /* (1, 26, 1) {real, imag} */,
  {32'hc438ac70, 32'h00000000} /* (1, 26, 0) {real, imag} */,
  {32'hc4d6fd9d, 32'h410ff680} /* (1, 25, 31) {real, imag} */,
  {32'h4419a775, 32'h42f9e4c5} /* (1, 25, 30) {real, imag} */,
  {32'h4101a8c7, 32'hc2831e7b} /* (1, 25, 29) {real, imag} */,
  {32'hc39ad8d3, 32'h426305e8} /* (1, 25, 28) {real, imag} */,
  {32'h431ba5ed, 32'hc2a21bc8} /* (1, 25, 27) {real, imag} */,
  {32'h428257a9, 32'hc1edd0d7} /* (1, 25, 26) {real, imag} */,
  {32'hc29f2eaf, 32'h432fa948} /* (1, 25, 25) {real, imag} */,
  {32'h40d522a0, 32'hc335205b} /* (1, 25, 24) {real, imag} */,
  {32'hc1a0c8a0, 32'hc249f2ce} /* (1, 25, 23) {real, imag} */,
  {32'hc227a526, 32'hc233e940} /* (1, 25, 22) {real, imag} */,
  {32'hc1971b00, 32'hc2e1d6d6} /* (1, 25, 21) {real, imag} */,
  {32'h420d9c9d, 32'hc2dcdc50} /* (1, 25, 20) {real, imag} */,
  {32'h42a56a03, 32'h4160f647} /* (1, 25, 19) {real, imag} */,
  {32'h40b57b44, 32'h415fddf4} /* (1, 25, 18) {real, imag} */,
  {32'h411a8c34, 32'hbfd155d8} /* (1, 25, 17) {real, imag} */,
  {32'h42a77bfb, 32'h00000000} /* (1, 25, 16) {real, imag} */,
  {32'h411a8c34, 32'h3fd155d8} /* (1, 25, 15) {real, imag} */,
  {32'h40b57b44, 32'hc15fddf4} /* (1, 25, 14) {real, imag} */,
  {32'h42a56a03, 32'hc160f647} /* (1, 25, 13) {real, imag} */,
  {32'h420d9c9d, 32'h42dcdc50} /* (1, 25, 12) {real, imag} */,
  {32'hc1971b00, 32'h42e1d6d6} /* (1, 25, 11) {real, imag} */,
  {32'hc227a526, 32'h4233e940} /* (1, 25, 10) {real, imag} */,
  {32'hc1a0c8a0, 32'h4249f2ce} /* (1, 25, 9) {real, imag} */,
  {32'h40d522a0, 32'h4335205b} /* (1, 25, 8) {real, imag} */,
  {32'hc29f2eaf, 32'hc32fa948} /* (1, 25, 7) {real, imag} */,
  {32'h428257a9, 32'h41edd0d7} /* (1, 25, 6) {real, imag} */,
  {32'h431ba5ed, 32'h42a21bc8} /* (1, 25, 5) {real, imag} */,
  {32'hc39ad8d3, 32'hc26305e8} /* (1, 25, 4) {real, imag} */,
  {32'h4101a8c7, 32'h42831e7b} /* (1, 25, 3) {real, imag} */,
  {32'h4419a775, 32'hc2f9e4c5} /* (1, 25, 2) {real, imag} */,
  {32'hc4d6fd9d, 32'hc10ff680} /* (1, 25, 1) {real, imag} */,
  {32'hc431851b, 32'h00000000} /* (1, 25, 0) {real, imag} */,
  {32'hc4c7d44c, 32'hc287782e} /* (1, 24, 31) {real, imag} */,
  {32'h4434db74, 32'h431c89ed} /* (1, 24, 30) {real, imag} */,
  {32'hc0f81630, 32'hc2979591} /* (1, 24, 29) {real, imag} */,
  {32'hc3a653a1, 32'hc191c83c} /* (1, 24, 28) {real, imag} */,
  {32'h435f35e2, 32'h40e0c080} /* (1, 24, 27) {real, imag} */,
  {32'hc218968c, 32'h417a5990} /* (1, 24, 26) {real, imag} */,
  {32'hc2377582, 32'h42d27f67} /* (1, 24, 25) {real, imag} */,
  {32'h424eb65a, 32'hc25abff7} /* (1, 24, 24) {real, imag} */,
  {32'h428619e0, 32'hc1b3fd08} /* (1, 24, 23) {real, imag} */,
  {32'hc23936d5, 32'h4298c915} /* (1, 24, 22) {real, imag} */,
  {32'h42897136, 32'hc29789d9} /* (1, 24, 21) {real, imag} */,
  {32'hc2b6b54a, 32'h42aaa458} /* (1, 24, 20) {real, imag} */,
  {32'h3f49b2e0, 32'h422db16a} /* (1, 24, 19) {real, imag} */,
  {32'h419e788a, 32'hc2b1fff0} /* (1, 24, 18) {real, imag} */,
  {32'hc200edb6, 32'h414f87a3} /* (1, 24, 17) {real, imag} */,
  {32'hc1960126, 32'h00000000} /* (1, 24, 16) {real, imag} */,
  {32'hc200edb6, 32'hc14f87a3} /* (1, 24, 15) {real, imag} */,
  {32'h419e788a, 32'h42b1fff0} /* (1, 24, 14) {real, imag} */,
  {32'h3f49b2e0, 32'hc22db16a} /* (1, 24, 13) {real, imag} */,
  {32'hc2b6b54a, 32'hc2aaa458} /* (1, 24, 12) {real, imag} */,
  {32'h42897136, 32'h429789d9} /* (1, 24, 11) {real, imag} */,
  {32'hc23936d5, 32'hc298c915} /* (1, 24, 10) {real, imag} */,
  {32'h428619e0, 32'h41b3fd08} /* (1, 24, 9) {real, imag} */,
  {32'h424eb65a, 32'h425abff7} /* (1, 24, 8) {real, imag} */,
  {32'hc2377582, 32'hc2d27f67} /* (1, 24, 7) {real, imag} */,
  {32'hc218968c, 32'hc17a5990} /* (1, 24, 6) {real, imag} */,
  {32'h435f35e2, 32'hc0e0c080} /* (1, 24, 5) {real, imag} */,
  {32'hc3a653a1, 32'h4191c83c} /* (1, 24, 4) {real, imag} */,
  {32'hc0f81630, 32'h42979591} /* (1, 24, 3) {real, imag} */,
  {32'h4434db74, 32'hc31c89ed} /* (1, 24, 2) {real, imag} */,
  {32'hc4c7d44c, 32'h4287782e} /* (1, 24, 1) {real, imag} */,
  {32'hc4030b24, 32'h00000000} /* (1, 24, 0) {real, imag} */,
  {32'hc4ae59d3, 32'h42473e7e} /* (1, 23, 31) {real, imag} */,
  {32'h43ecad30, 32'h42b3e9f1} /* (1, 23, 30) {real, imag} */,
  {32'h42cac1c8, 32'h41cf6dc6} /* (1, 23, 29) {real, imag} */,
  {32'hc377f5ae, 32'h40afe114} /* (1, 23, 28) {real, imag} */,
  {32'h428370d5, 32'hc2e7fb71} /* (1, 23, 27) {real, imag} */,
  {32'h42237838, 32'h42695115} /* (1, 23, 26) {real, imag} */,
  {32'hc1da04cc, 32'h428bf520} /* (1, 23, 25) {real, imag} */,
  {32'h41423270, 32'hc2936ce2} /* (1, 23, 24) {real, imag} */,
  {32'h41890571, 32'hc25f2e9c} /* (1, 23, 23) {real, imag} */,
  {32'h41ec3781, 32'hc232fac7} /* (1, 23, 22) {real, imag} */,
  {32'h4239c8f5, 32'hc285fa54} /* (1, 23, 21) {real, imag} */,
  {32'h41df917c, 32'h426ccb33} /* (1, 23, 20) {real, imag} */,
  {32'hc138578e, 32'h41dff9c6} /* (1, 23, 19) {real, imag} */,
  {32'h420ad3b6, 32'hc2cb671e} /* (1, 23, 18) {real, imag} */,
  {32'h425411d3, 32'h42b54013} /* (1, 23, 17) {real, imag} */,
  {32'h40ed7046, 32'h00000000} /* (1, 23, 16) {real, imag} */,
  {32'h425411d3, 32'hc2b54013} /* (1, 23, 15) {real, imag} */,
  {32'h420ad3b6, 32'h42cb671e} /* (1, 23, 14) {real, imag} */,
  {32'hc138578e, 32'hc1dff9c6} /* (1, 23, 13) {real, imag} */,
  {32'h41df917c, 32'hc26ccb33} /* (1, 23, 12) {real, imag} */,
  {32'h4239c8f5, 32'h4285fa54} /* (1, 23, 11) {real, imag} */,
  {32'h41ec3781, 32'h4232fac7} /* (1, 23, 10) {real, imag} */,
  {32'h41890571, 32'h425f2e9c} /* (1, 23, 9) {real, imag} */,
  {32'h41423270, 32'h42936ce2} /* (1, 23, 8) {real, imag} */,
  {32'hc1da04cc, 32'hc28bf520} /* (1, 23, 7) {real, imag} */,
  {32'h42237838, 32'hc2695115} /* (1, 23, 6) {real, imag} */,
  {32'h428370d5, 32'h42e7fb71} /* (1, 23, 5) {real, imag} */,
  {32'hc377f5ae, 32'hc0afe114} /* (1, 23, 4) {real, imag} */,
  {32'h42cac1c8, 32'hc1cf6dc6} /* (1, 23, 3) {real, imag} */,
  {32'h43ecad30, 32'hc2b3e9f1} /* (1, 23, 2) {real, imag} */,
  {32'hc4ae59d3, 32'hc2473e7e} /* (1, 23, 1) {real, imag} */,
  {32'hc39f8856, 32'h00000000} /* (1, 23, 0) {real, imag} */,
  {32'hc48a61c2, 32'h42ae4d6e} /* (1, 22, 31) {real, imag} */,
  {32'h43dadfde, 32'h428bee02} /* (1, 22, 30) {real, imag} */,
  {32'h42d639c5, 32'h429ecac8} /* (1, 22, 29) {real, imag} */,
  {32'hc2ff5d78, 32'hc2c2daf8} /* (1, 22, 28) {real, imag} */,
  {32'h42a3b576, 32'hc330f0b0} /* (1, 22, 27) {real, imag} */,
  {32'hc222ddea, 32'h40a330f6} /* (1, 22, 26) {real, imag} */,
  {32'hc31348b4, 32'h427ffc2b} /* (1, 22, 25) {real, imag} */,
  {32'h4265d528, 32'hc21a6e71} /* (1, 22, 24) {real, imag} */,
  {32'hc28e4f60, 32'h41bccd2d} /* (1, 22, 23) {real, imag} */,
  {32'h42bd85ad, 32'h430d8bb4} /* (1, 22, 22) {real, imag} */,
  {32'h41dc4ebe, 32'hc25afe8a} /* (1, 22, 21) {real, imag} */,
  {32'h41d087d1, 32'h42065f5c} /* (1, 22, 20) {real, imag} */,
  {32'h4186f24b, 32'hc134d51c} /* (1, 22, 19) {real, imag} */,
  {32'h416df7e0, 32'hc1c9ba6c} /* (1, 22, 18) {real, imag} */,
  {32'hc1d087f1, 32'h4190c1be} /* (1, 22, 17) {real, imag} */,
  {32'h42a0bf8e, 32'h00000000} /* (1, 22, 16) {real, imag} */,
  {32'hc1d087f1, 32'hc190c1be} /* (1, 22, 15) {real, imag} */,
  {32'h416df7e0, 32'h41c9ba6c} /* (1, 22, 14) {real, imag} */,
  {32'h4186f24b, 32'h4134d51c} /* (1, 22, 13) {real, imag} */,
  {32'h41d087d1, 32'hc2065f5c} /* (1, 22, 12) {real, imag} */,
  {32'h41dc4ebe, 32'h425afe8a} /* (1, 22, 11) {real, imag} */,
  {32'h42bd85ad, 32'hc30d8bb4} /* (1, 22, 10) {real, imag} */,
  {32'hc28e4f60, 32'hc1bccd2d} /* (1, 22, 9) {real, imag} */,
  {32'h4265d528, 32'h421a6e71} /* (1, 22, 8) {real, imag} */,
  {32'hc31348b4, 32'hc27ffc2b} /* (1, 22, 7) {real, imag} */,
  {32'hc222ddea, 32'hc0a330f6} /* (1, 22, 6) {real, imag} */,
  {32'h42a3b576, 32'h4330f0b0} /* (1, 22, 5) {real, imag} */,
  {32'hc2ff5d78, 32'h42c2daf8} /* (1, 22, 4) {real, imag} */,
  {32'h42d639c5, 32'hc29ecac8} /* (1, 22, 3) {real, imag} */,
  {32'h43dadfde, 32'hc28bee02} /* (1, 22, 2) {real, imag} */,
  {32'hc48a61c2, 32'hc2ae4d6e} /* (1, 22, 1) {real, imag} */,
  {32'hc3600bf6, 32'h00000000} /* (1, 22, 0) {real, imag} */,
  {32'hc3e6dfd4, 32'h41933588} /* (1, 21, 31) {real, imag} */,
  {32'h4300e04c, 32'h40833600} /* (1, 21, 30) {real, imag} */,
  {32'hc1b1a0b7, 32'h42f0397b} /* (1, 21, 29) {real, imag} */,
  {32'hc2d19bd6, 32'h41a06bc0} /* (1, 21, 28) {real, imag} */,
  {32'h4262ec50, 32'hc261b87f} /* (1, 21, 27) {real, imag} */,
  {32'hc24200a8, 32'h3f8cf040} /* (1, 21, 26) {real, imag} */,
  {32'hc223742d, 32'h4250f97e} /* (1, 21, 25) {real, imag} */,
  {32'hc29e1288, 32'hc20f3287} /* (1, 21, 24) {real, imag} */,
  {32'h424b1d70, 32'h42cc97ac} /* (1, 21, 23) {real, imag} */,
  {32'h425602e4, 32'h41cd8904} /* (1, 21, 22) {real, imag} */,
  {32'h42a2813e, 32'h42adfcc7} /* (1, 21, 21) {real, imag} */,
  {32'h4267b6ad, 32'hc2676b67} /* (1, 21, 20) {real, imag} */,
  {32'h423bea8a, 32'h41b969e8} /* (1, 21, 19) {real, imag} */,
  {32'h41215b2f, 32'hc2217a5f} /* (1, 21, 18) {real, imag} */,
  {32'hc1dfd983, 32'hc0e0297c} /* (1, 21, 17) {real, imag} */,
  {32'hc25c51b7, 32'h00000000} /* (1, 21, 16) {real, imag} */,
  {32'hc1dfd983, 32'h40e0297c} /* (1, 21, 15) {real, imag} */,
  {32'h41215b2f, 32'h42217a5f} /* (1, 21, 14) {real, imag} */,
  {32'h423bea8a, 32'hc1b969e8} /* (1, 21, 13) {real, imag} */,
  {32'h4267b6ad, 32'h42676b67} /* (1, 21, 12) {real, imag} */,
  {32'h42a2813e, 32'hc2adfcc7} /* (1, 21, 11) {real, imag} */,
  {32'h425602e4, 32'hc1cd8904} /* (1, 21, 10) {real, imag} */,
  {32'h424b1d70, 32'hc2cc97ac} /* (1, 21, 9) {real, imag} */,
  {32'hc29e1288, 32'h420f3287} /* (1, 21, 8) {real, imag} */,
  {32'hc223742d, 32'hc250f97e} /* (1, 21, 7) {real, imag} */,
  {32'hc24200a8, 32'hbf8cf040} /* (1, 21, 6) {real, imag} */,
  {32'h4262ec50, 32'h4261b87f} /* (1, 21, 5) {real, imag} */,
  {32'hc2d19bd6, 32'hc1a06bc0} /* (1, 21, 4) {real, imag} */,
  {32'hc1b1a0b7, 32'hc2f0397b} /* (1, 21, 3) {real, imag} */,
  {32'h4300e04c, 32'hc0833600} /* (1, 21, 2) {real, imag} */,
  {32'hc3e6dfd4, 32'hc1933588} /* (1, 21, 1) {real, imag} */,
  {32'hc1ce0f30, 32'h00000000} /* (1, 21, 0) {real, imag} */,
  {32'h440e253e, 32'hc37f4662} /* (1, 20, 31) {real, imag} */,
  {32'hc3d3f884, 32'h4254f71f} /* (1, 20, 30) {real, imag} */,
  {32'h420a913c, 32'h43097154} /* (1, 20, 29) {real, imag} */,
  {32'hc10f99a0, 32'hc2873e53} /* (1, 20, 28) {real, imag} */,
  {32'hc300d642, 32'h41fd5a2c} /* (1, 20, 27) {real, imag} */,
  {32'hc2e54076, 32'h426ba22b} /* (1, 20, 26) {real, imag} */,
  {32'hc2b228d0, 32'h3f673f10} /* (1, 20, 25) {real, imag} */,
  {32'hc25524c8, 32'h42ec63b1} /* (1, 20, 24) {real, imag} */,
  {32'h417f6824, 32'hc2a5349c} /* (1, 20, 23) {real, imag} */,
  {32'hc19961c2, 32'hc2637b65} /* (1, 20, 22) {real, imag} */,
  {32'hc278cad8, 32'hc28b2442} /* (1, 20, 21) {real, imag} */,
  {32'hc1988273, 32'h425f0aa6} /* (1, 20, 20) {real, imag} */,
  {32'h41d0f7e2, 32'hc285d476} /* (1, 20, 19) {real, imag} */,
  {32'h41913bb8, 32'hc24b843c} /* (1, 20, 18) {real, imag} */,
  {32'hc20a25f1, 32'hc1af65bc} /* (1, 20, 17) {real, imag} */,
  {32'h41c59bce, 32'h00000000} /* (1, 20, 16) {real, imag} */,
  {32'hc20a25f1, 32'h41af65bc} /* (1, 20, 15) {real, imag} */,
  {32'h41913bb8, 32'h424b843c} /* (1, 20, 14) {real, imag} */,
  {32'h41d0f7e2, 32'h4285d476} /* (1, 20, 13) {real, imag} */,
  {32'hc1988273, 32'hc25f0aa6} /* (1, 20, 12) {real, imag} */,
  {32'hc278cad8, 32'h428b2442} /* (1, 20, 11) {real, imag} */,
  {32'hc19961c2, 32'h42637b65} /* (1, 20, 10) {real, imag} */,
  {32'h417f6824, 32'h42a5349c} /* (1, 20, 9) {real, imag} */,
  {32'hc25524c8, 32'hc2ec63b1} /* (1, 20, 8) {real, imag} */,
  {32'hc2b228d0, 32'hbf673f10} /* (1, 20, 7) {real, imag} */,
  {32'hc2e54076, 32'hc26ba22b} /* (1, 20, 6) {real, imag} */,
  {32'hc300d642, 32'hc1fd5a2c} /* (1, 20, 5) {real, imag} */,
  {32'hc10f99a0, 32'h42873e53} /* (1, 20, 4) {real, imag} */,
  {32'h420a913c, 32'hc3097154} /* (1, 20, 3) {real, imag} */,
  {32'hc3d3f884, 32'hc254f71f} /* (1, 20, 2) {real, imag} */,
  {32'h440e253e, 32'h437f4662} /* (1, 20, 1) {real, imag} */,
  {32'h44111036, 32'h00000000} /* (1, 20, 0) {real, imag} */,
  {32'h44836bc5, 32'hc39a26bc} /* (1, 19, 31) {real, imag} */,
  {32'hc40ff06a, 32'h437f9082} /* (1, 19, 30) {real, imag} */,
  {32'hc0c81d08, 32'h43035c07} /* (1, 19, 29) {real, imag} */,
  {32'h42e818a7, 32'hc31a54e0} /* (1, 19, 28) {real, imag} */,
  {32'hc31453e6, 32'h426cbe24} /* (1, 19, 27) {real, imag} */,
  {32'hc268768f, 32'hc1ca4963} /* (1, 19, 26) {real, imag} */,
  {32'h41b167b3, 32'hc28d828a} /* (1, 19, 25) {real, imag} */,
  {32'hc20ebebd, 32'hc172b4dc} /* (1, 19, 24) {real, imag} */,
  {32'h423de9b4, 32'h41aa027e} /* (1, 19, 23) {real, imag} */,
  {32'h4236de56, 32'h418cc30f} /* (1, 19, 22) {real, imag} */,
  {32'hc1a8677e, 32'h42034898} /* (1, 19, 21) {real, imag} */,
  {32'h41628404, 32'h4278e4fa} /* (1, 19, 20) {real, imag} */,
  {32'hc17989e8, 32'h4230e8d2} /* (1, 19, 19) {real, imag} */,
  {32'hc1857b5d, 32'h41dbe43e} /* (1, 19, 18) {real, imag} */,
  {32'hc2363627, 32'hc206380e} /* (1, 19, 17) {real, imag} */,
  {32'hc31902e2, 32'h00000000} /* (1, 19, 16) {real, imag} */,
  {32'hc2363627, 32'h4206380e} /* (1, 19, 15) {real, imag} */,
  {32'hc1857b5d, 32'hc1dbe43e} /* (1, 19, 14) {real, imag} */,
  {32'hc17989e8, 32'hc230e8d2} /* (1, 19, 13) {real, imag} */,
  {32'h41628404, 32'hc278e4fa} /* (1, 19, 12) {real, imag} */,
  {32'hc1a8677e, 32'hc2034898} /* (1, 19, 11) {real, imag} */,
  {32'h4236de56, 32'hc18cc30f} /* (1, 19, 10) {real, imag} */,
  {32'h423de9b4, 32'hc1aa027e} /* (1, 19, 9) {real, imag} */,
  {32'hc20ebebd, 32'h4172b4dc} /* (1, 19, 8) {real, imag} */,
  {32'h41b167b3, 32'h428d828a} /* (1, 19, 7) {real, imag} */,
  {32'hc268768f, 32'h41ca4963} /* (1, 19, 6) {real, imag} */,
  {32'hc31453e6, 32'hc26cbe24} /* (1, 19, 5) {real, imag} */,
  {32'h42e818a7, 32'h431a54e0} /* (1, 19, 4) {real, imag} */,
  {32'hc0c81d08, 32'hc3035c07} /* (1, 19, 3) {real, imag} */,
  {32'hc40ff06a, 32'hc37f9082} /* (1, 19, 2) {real, imag} */,
  {32'h44836bc5, 32'h439a26bc} /* (1, 19, 1) {real, imag} */,
  {32'h446f3bd3, 32'h00000000} /* (1, 19, 0) {real, imag} */,
  {32'h448fe388, 32'hc353e288} /* (1, 18, 31) {real, imag} */,
  {32'hc4342999, 32'h43005f76} /* (1, 18, 30) {real, imag} */,
  {32'hc257d53e, 32'h419a54af} /* (1, 18, 29) {real, imag} */,
  {32'h43429720, 32'h41bdc0d6} /* (1, 18, 28) {real, imag} */,
  {32'hc2b5ef13, 32'h4239919f} /* (1, 18, 27) {real, imag} */,
  {32'h4241d45c, 32'h40324f90} /* (1, 18, 26) {real, imag} */,
  {32'hc20b69d5, 32'hc24ce911} /* (1, 18, 25) {real, imag} */,
  {32'hc28e58d0, 32'hc30697f7} /* (1, 18, 24) {real, imag} */,
  {32'hc10cbeb0, 32'h41c97012} /* (1, 18, 23) {real, imag} */,
  {32'h4206ec3a, 32'h419c1ccf} /* (1, 18, 22) {real, imag} */,
  {32'hc07f9bf8, 32'h427ae7fe} /* (1, 18, 21) {real, imag} */,
  {32'h410d1fae, 32'hc221ebac} /* (1, 18, 20) {real, imag} */,
  {32'h430ef2a9, 32'hc295fc0c} /* (1, 18, 19) {real, imag} */,
  {32'h429ce1d4, 32'h41e682e4} /* (1, 18, 18) {real, imag} */,
  {32'h4178335c, 32'h428add3c} /* (1, 18, 17) {real, imag} */,
  {32'h42568417, 32'h00000000} /* (1, 18, 16) {real, imag} */,
  {32'h4178335c, 32'hc28add3c} /* (1, 18, 15) {real, imag} */,
  {32'h429ce1d4, 32'hc1e682e4} /* (1, 18, 14) {real, imag} */,
  {32'h430ef2a9, 32'h4295fc0c} /* (1, 18, 13) {real, imag} */,
  {32'h410d1fae, 32'h4221ebac} /* (1, 18, 12) {real, imag} */,
  {32'hc07f9bf8, 32'hc27ae7fe} /* (1, 18, 11) {real, imag} */,
  {32'h4206ec3a, 32'hc19c1ccf} /* (1, 18, 10) {real, imag} */,
  {32'hc10cbeb0, 32'hc1c97012} /* (1, 18, 9) {real, imag} */,
  {32'hc28e58d0, 32'h430697f7} /* (1, 18, 8) {real, imag} */,
  {32'hc20b69d5, 32'h424ce911} /* (1, 18, 7) {real, imag} */,
  {32'h4241d45c, 32'hc0324f90} /* (1, 18, 6) {real, imag} */,
  {32'hc2b5ef13, 32'hc239919f} /* (1, 18, 5) {real, imag} */,
  {32'h43429720, 32'hc1bdc0d6} /* (1, 18, 4) {real, imag} */,
  {32'hc257d53e, 32'hc19a54af} /* (1, 18, 3) {real, imag} */,
  {32'hc4342999, 32'hc3005f76} /* (1, 18, 2) {real, imag} */,
  {32'h448fe388, 32'h4353e288} /* (1, 18, 1) {real, imag} */,
  {32'h4482a12b, 32'h00000000} /* (1, 18, 0) {real, imag} */,
  {32'h44a434e2, 32'hc3802c4b} /* (1, 17, 31) {real, imag} */,
  {32'hc454b398, 32'h425b086c} /* (1, 17, 30) {real, imag} */,
  {32'hc223422d, 32'hc283d1ed} /* (1, 17, 29) {real, imag} */,
  {32'h43415f48, 32'hc301e2b4} /* (1, 17, 28) {real, imag} */,
  {32'hc2c15ba3, 32'h425f9782} /* (1, 17, 27) {real, imag} */,
  {32'h42280145, 32'hc1f1daac} /* (1, 17, 26) {real, imag} */,
  {32'h42d8c955, 32'h41b90418} /* (1, 17, 25) {real, imag} */,
  {32'hc3291aae, 32'hbeeba000} /* (1, 17, 24) {real, imag} */,
  {32'hc28d2327, 32'hc166bfe8} /* (1, 17, 23) {real, imag} */,
  {32'h42050a41, 32'hc258189e} /* (1, 17, 22) {real, imag} */,
  {32'hc05a46c8, 32'hc29fc8ec} /* (1, 17, 21) {real, imag} */,
  {32'hc2a96cf2, 32'h42d34791} /* (1, 17, 20) {real, imag} */,
  {32'h40c548e0, 32'h42ba4be9} /* (1, 17, 19) {real, imag} */,
  {32'hc23475fa, 32'hc16c0aef} /* (1, 17, 18) {real, imag} */,
  {32'hc1a61bae, 32'hc2854aeb} /* (1, 17, 17) {real, imag} */,
  {32'h42a12d8d, 32'h00000000} /* (1, 17, 16) {real, imag} */,
  {32'hc1a61bae, 32'h42854aeb} /* (1, 17, 15) {real, imag} */,
  {32'hc23475fa, 32'h416c0aef} /* (1, 17, 14) {real, imag} */,
  {32'h40c548e0, 32'hc2ba4be9} /* (1, 17, 13) {real, imag} */,
  {32'hc2a96cf2, 32'hc2d34791} /* (1, 17, 12) {real, imag} */,
  {32'hc05a46c8, 32'h429fc8ec} /* (1, 17, 11) {real, imag} */,
  {32'h42050a41, 32'h4258189e} /* (1, 17, 10) {real, imag} */,
  {32'hc28d2327, 32'h4166bfe8} /* (1, 17, 9) {real, imag} */,
  {32'hc3291aae, 32'h3eeba000} /* (1, 17, 8) {real, imag} */,
  {32'h42d8c955, 32'hc1b90418} /* (1, 17, 7) {real, imag} */,
  {32'h42280145, 32'h41f1daac} /* (1, 17, 6) {real, imag} */,
  {32'hc2c15ba3, 32'hc25f9782} /* (1, 17, 5) {real, imag} */,
  {32'h43415f48, 32'h4301e2b4} /* (1, 17, 4) {real, imag} */,
  {32'hc223422d, 32'h4283d1ed} /* (1, 17, 3) {real, imag} */,
  {32'hc454b398, 32'hc25b086c} /* (1, 17, 2) {real, imag} */,
  {32'h44a434e2, 32'h43802c4b} /* (1, 17, 1) {real, imag} */,
  {32'h44934e21, 32'h00000000} /* (1, 17, 0) {real, imag} */,
  {32'h44aa108c, 32'hc364ace8} /* (1, 16, 31) {real, imag} */,
  {32'hc4546434, 32'h42f37dc4} /* (1, 16, 30) {real, imag} */,
  {32'h428bb28e, 32'hc302ba4b} /* (1, 16, 29) {real, imag} */,
  {32'h4317fee8, 32'hc30bfb73} /* (1, 16, 28) {real, imag} */,
  {32'hc2c3b84e, 32'h434fec0c} /* (1, 16, 27) {real, imag} */,
  {32'h428a3583, 32'h42863507} /* (1, 16, 26) {real, imag} */,
  {32'h4292639c, 32'hc1cc4d6a} /* (1, 16, 25) {real, imag} */,
  {32'hc29c1be8, 32'h4301831e} /* (1, 16, 24) {real, imag} */,
  {32'hbf2b26c0, 32'h4256aa1d} /* (1, 16, 23) {real, imag} */,
  {32'h42cc64f6, 32'hc265d2ef} /* (1, 16, 22) {real, imag} */,
  {32'h41018bba, 32'h42984e96} /* (1, 16, 21) {real, imag} */,
  {32'hc1b02530, 32'h42850c8f} /* (1, 16, 20) {real, imag} */,
  {32'hc1bb0266, 32'h41f934de} /* (1, 16, 19) {real, imag} */,
  {32'h41f20280, 32'hc204e9ac} /* (1, 16, 18) {real, imag} */,
  {32'hc0f5a8de, 32'hc17173db} /* (1, 16, 17) {real, imag} */,
  {32'hc2219806, 32'h00000000} /* (1, 16, 16) {real, imag} */,
  {32'hc0f5a8de, 32'h417173db} /* (1, 16, 15) {real, imag} */,
  {32'h41f20280, 32'h4204e9ac} /* (1, 16, 14) {real, imag} */,
  {32'hc1bb0266, 32'hc1f934de} /* (1, 16, 13) {real, imag} */,
  {32'hc1b02530, 32'hc2850c8f} /* (1, 16, 12) {real, imag} */,
  {32'h41018bba, 32'hc2984e96} /* (1, 16, 11) {real, imag} */,
  {32'h42cc64f6, 32'h4265d2ef} /* (1, 16, 10) {real, imag} */,
  {32'hbf2b26c0, 32'hc256aa1d} /* (1, 16, 9) {real, imag} */,
  {32'hc29c1be8, 32'hc301831e} /* (1, 16, 8) {real, imag} */,
  {32'h4292639c, 32'h41cc4d6a} /* (1, 16, 7) {real, imag} */,
  {32'h428a3583, 32'hc2863507} /* (1, 16, 6) {real, imag} */,
  {32'hc2c3b84e, 32'hc34fec0c} /* (1, 16, 5) {real, imag} */,
  {32'h4317fee8, 32'h430bfb73} /* (1, 16, 4) {real, imag} */,
  {32'h428bb28e, 32'h4302ba4b} /* (1, 16, 3) {real, imag} */,
  {32'hc4546434, 32'hc2f37dc4} /* (1, 16, 2) {real, imag} */,
  {32'h44aa108c, 32'h4364ace8} /* (1, 16, 1) {real, imag} */,
  {32'h448c1a27, 32'h00000000} /* (1, 16, 0) {real, imag} */,
  {32'h44c2f082, 32'hc35ad89a} /* (1, 15, 31) {real, imag} */,
  {32'hc426349c, 32'h432fcbe5} /* (1, 15, 30) {real, imag} */,
  {32'hc28e058a, 32'hc2ad3069} /* (1, 15, 29) {real, imag} */,
  {32'h430a64b0, 32'hc2a281a1} /* (1, 15, 28) {real, imag} */,
  {32'hc32d4514, 32'h4321aaac} /* (1, 15, 27) {real, imag} */,
  {32'h41d7d1ea, 32'h425c5072} /* (1, 15, 26) {real, imag} */,
  {32'h41bab43c, 32'h4139e9a4} /* (1, 15, 25) {real, imag} */,
  {32'hc2d31243, 32'h4313f86c} /* (1, 15, 24) {real, imag} */,
  {32'h42ba7ae5, 32'h425679b6} /* (1, 15, 23) {real, imag} */,
  {32'hc24d8c7d, 32'h4190a11f} /* (1, 15, 22) {real, imag} */,
  {32'h41bce23d, 32'h42bf9e44} /* (1, 15, 21) {real, imag} */,
  {32'hc1bb82ee, 32'h41204aa8} /* (1, 15, 20) {real, imag} */,
  {32'hc25324f2, 32'hc297d233} /* (1, 15, 19) {real, imag} */,
  {32'hc2221516, 32'hc1a3293a} /* (1, 15, 18) {real, imag} */,
  {32'h416f8974, 32'hc0f0c634} /* (1, 15, 17) {real, imag} */,
  {32'hc21db93a, 32'h00000000} /* (1, 15, 16) {real, imag} */,
  {32'h416f8974, 32'h40f0c634} /* (1, 15, 15) {real, imag} */,
  {32'hc2221516, 32'h41a3293a} /* (1, 15, 14) {real, imag} */,
  {32'hc25324f2, 32'h4297d233} /* (1, 15, 13) {real, imag} */,
  {32'hc1bb82ee, 32'hc1204aa8} /* (1, 15, 12) {real, imag} */,
  {32'h41bce23d, 32'hc2bf9e44} /* (1, 15, 11) {real, imag} */,
  {32'hc24d8c7d, 32'hc190a11f} /* (1, 15, 10) {real, imag} */,
  {32'h42ba7ae5, 32'hc25679b6} /* (1, 15, 9) {real, imag} */,
  {32'hc2d31243, 32'hc313f86c} /* (1, 15, 8) {real, imag} */,
  {32'h41bab43c, 32'hc139e9a4} /* (1, 15, 7) {real, imag} */,
  {32'h41d7d1ea, 32'hc25c5072} /* (1, 15, 6) {real, imag} */,
  {32'hc32d4514, 32'hc321aaac} /* (1, 15, 5) {real, imag} */,
  {32'h430a64b0, 32'h42a281a1} /* (1, 15, 4) {real, imag} */,
  {32'hc28e058a, 32'h42ad3069} /* (1, 15, 3) {real, imag} */,
  {32'hc426349c, 32'hc32fcbe5} /* (1, 15, 2) {real, imag} */,
  {32'h44c2f082, 32'h435ad89a} /* (1, 15, 1) {real, imag} */,
  {32'h448e3dc1, 32'h00000000} /* (1, 15, 0) {real, imag} */,
  {32'h44d10e34, 32'hc38a0872} /* (1, 14, 31) {real, imag} */,
  {32'hc433b965, 32'h4297c60c} /* (1, 14, 30) {real, imag} */,
  {32'hc2226d0a, 32'hc27f401c} /* (1, 14, 29) {real, imag} */,
  {32'h42e3b0f7, 32'hc2878ea4} /* (1, 14, 28) {real, imag} */,
  {32'hc3771f06, 32'h42e2d778} /* (1, 14, 27) {real, imag} */,
  {32'h42418064, 32'hc29f894c} /* (1, 14, 26) {real, imag} */,
  {32'hc2b427cc, 32'h3e7f2500} /* (1, 14, 25) {real, imag} */,
  {32'hc298d844, 32'hc16e7494} /* (1, 14, 24) {real, imag} */,
  {32'hc2b56556, 32'h42684687} /* (1, 14, 23) {real, imag} */,
  {32'h40b9cfc0, 32'hc0c02c94} /* (1, 14, 22) {real, imag} */,
  {32'hc268b4dc, 32'h41d5c018} /* (1, 14, 21) {real, imag} */,
  {32'h424f7d5e, 32'h421ff73e} /* (1, 14, 20) {real, imag} */,
  {32'hc1750990, 32'h40cbc600} /* (1, 14, 19) {real, imag} */,
  {32'h41a983f6, 32'h411065e0} /* (1, 14, 18) {real, imag} */,
  {32'hc29659b8, 32'hc0bb2ec0} /* (1, 14, 17) {real, imag} */,
  {32'h42bd908c, 32'h00000000} /* (1, 14, 16) {real, imag} */,
  {32'hc29659b8, 32'h40bb2ec0} /* (1, 14, 15) {real, imag} */,
  {32'h41a983f6, 32'hc11065e0} /* (1, 14, 14) {real, imag} */,
  {32'hc1750990, 32'hc0cbc600} /* (1, 14, 13) {real, imag} */,
  {32'h424f7d5e, 32'hc21ff73e} /* (1, 14, 12) {real, imag} */,
  {32'hc268b4dc, 32'hc1d5c018} /* (1, 14, 11) {real, imag} */,
  {32'h40b9cfc0, 32'h40c02c94} /* (1, 14, 10) {real, imag} */,
  {32'hc2b56556, 32'hc2684687} /* (1, 14, 9) {real, imag} */,
  {32'hc298d844, 32'h416e7494} /* (1, 14, 8) {real, imag} */,
  {32'hc2b427cc, 32'hbe7f2500} /* (1, 14, 7) {real, imag} */,
  {32'h42418064, 32'h429f894c} /* (1, 14, 6) {real, imag} */,
  {32'hc3771f06, 32'hc2e2d778} /* (1, 14, 5) {real, imag} */,
  {32'h42e3b0f7, 32'h42878ea4} /* (1, 14, 4) {real, imag} */,
  {32'hc2226d0a, 32'h427f401c} /* (1, 14, 3) {real, imag} */,
  {32'hc433b965, 32'hc297c60c} /* (1, 14, 2) {real, imag} */,
  {32'h44d10e34, 32'h438a0872} /* (1, 14, 1) {real, imag} */,
  {32'h4476427b, 32'h00000000} /* (1, 14, 0) {real, imag} */,
  {32'h44cf8c97, 32'hc38e6f30} /* (1, 13, 31) {real, imag} */,
  {32'hc4390aa6, 32'hc21b1cc0} /* (1, 13, 30) {real, imag} */,
  {32'hc234ee3d, 32'h41fe7df8} /* (1, 13, 29) {real, imag} */,
  {32'h42b77749, 32'hc2a41721} /* (1, 13, 28) {real, imag} */,
  {32'hc2e9130f, 32'h4394af30} /* (1, 13, 27) {real, imag} */,
  {32'hc2cadbfe, 32'hc1f36c99} /* (1, 13, 26) {real, imag} */,
  {32'h41cdf32d, 32'hc28c258c} /* (1, 13, 25) {real, imag} */,
  {32'hc2bd3be2, 32'h42cab50e} /* (1, 13, 24) {real, imag} */,
  {32'h426bc4ba, 32'h429d3a40} /* (1, 13, 23) {real, imag} */,
  {32'hc1f4f6c4, 32'hc1be4c41} /* (1, 13, 22) {real, imag} */,
  {32'h4238fd05, 32'hc1fecea8} /* (1, 13, 21) {real, imag} */,
  {32'h41b79ad2, 32'hc2f3b1dd} /* (1, 13, 20) {real, imag} */,
  {32'h431cd578, 32'hc11f0466} /* (1, 13, 19) {real, imag} */,
  {32'hc11657fe, 32'hc21598a9} /* (1, 13, 18) {real, imag} */,
  {32'h3fed0260, 32'h411e3d8e} /* (1, 13, 17) {real, imag} */,
  {32'hc1e57d50, 32'h00000000} /* (1, 13, 16) {real, imag} */,
  {32'h3fed0260, 32'hc11e3d8e} /* (1, 13, 15) {real, imag} */,
  {32'hc11657fe, 32'h421598a9} /* (1, 13, 14) {real, imag} */,
  {32'h431cd578, 32'h411f0466} /* (1, 13, 13) {real, imag} */,
  {32'h41b79ad2, 32'h42f3b1dd} /* (1, 13, 12) {real, imag} */,
  {32'h4238fd05, 32'h41fecea8} /* (1, 13, 11) {real, imag} */,
  {32'hc1f4f6c4, 32'h41be4c41} /* (1, 13, 10) {real, imag} */,
  {32'h426bc4ba, 32'hc29d3a40} /* (1, 13, 9) {real, imag} */,
  {32'hc2bd3be2, 32'hc2cab50e} /* (1, 13, 8) {real, imag} */,
  {32'h41cdf32d, 32'h428c258c} /* (1, 13, 7) {real, imag} */,
  {32'hc2cadbfe, 32'h41f36c99} /* (1, 13, 6) {real, imag} */,
  {32'hc2e9130f, 32'hc394af30} /* (1, 13, 5) {real, imag} */,
  {32'h42b77749, 32'h42a41721} /* (1, 13, 4) {real, imag} */,
  {32'hc234ee3d, 32'hc1fe7df8} /* (1, 13, 3) {real, imag} */,
  {32'hc4390aa6, 32'h421b1cc0} /* (1, 13, 2) {real, imag} */,
  {32'h44cf8c97, 32'h438e6f30} /* (1, 13, 1) {real, imag} */,
  {32'h445b1b69, 32'h00000000} /* (1, 13, 0) {real, imag} */,
  {32'h44a5c934, 32'hc381e1f3} /* (1, 12, 31) {real, imag} */,
  {32'hc42fd606, 32'h42beda28} /* (1, 12, 30) {real, imag} */,
  {32'h41c93e6c, 32'h43210d70} /* (1, 12, 29) {real, imag} */,
  {32'h42eb9b40, 32'hc35fcfe4} /* (1, 12, 28) {real, imag} */,
  {32'hc32b5470, 32'h431258f2} /* (1, 12, 27) {real, imag} */,
  {32'hc20e38a4, 32'h4292fadf} /* (1, 12, 26) {real, imag} */,
  {32'h4321aa2a, 32'h41934ef8} /* (1, 12, 25) {real, imag} */,
  {32'hc28ef25b, 32'h4216fb46} /* (1, 12, 24) {real, imag} */,
  {32'h41f69656, 32'h40658e10} /* (1, 12, 23) {real, imag} */,
  {32'h419ed070, 32'hc1c9b2de} /* (1, 12, 22) {real, imag} */,
  {32'h429a11b0, 32'h4301b501} /* (1, 12, 21) {real, imag} */,
  {32'hc2010f75, 32'hc2c1583d} /* (1, 12, 20) {real, imag} */,
  {32'h41b0dda2, 32'h425e18a9} /* (1, 12, 19) {real, imag} */,
  {32'h40e18860, 32'h424156cc} /* (1, 12, 18) {real, imag} */,
  {32'hc1869086, 32'h41bf94f0} /* (1, 12, 17) {real, imag} */,
  {32'h41ad50f8, 32'h00000000} /* (1, 12, 16) {real, imag} */,
  {32'hc1869086, 32'hc1bf94f0} /* (1, 12, 15) {real, imag} */,
  {32'h40e18860, 32'hc24156cc} /* (1, 12, 14) {real, imag} */,
  {32'h41b0dda2, 32'hc25e18a9} /* (1, 12, 13) {real, imag} */,
  {32'hc2010f75, 32'h42c1583d} /* (1, 12, 12) {real, imag} */,
  {32'h429a11b0, 32'hc301b501} /* (1, 12, 11) {real, imag} */,
  {32'h419ed070, 32'h41c9b2de} /* (1, 12, 10) {real, imag} */,
  {32'h41f69656, 32'hc0658e10} /* (1, 12, 9) {real, imag} */,
  {32'hc28ef25b, 32'hc216fb46} /* (1, 12, 8) {real, imag} */,
  {32'h4321aa2a, 32'hc1934ef8} /* (1, 12, 7) {real, imag} */,
  {32'hc20e38a4, 32'hc292fadf} /* (1, 12, 6) {real, imag} */,
  {32'hc32b5470, 32'hc31258f2} /* (1, 12, 5) {real, imag} */,
  {32'h42eb9b40, 32'h435fcfe4} /* (1, 12, 4) {real, imag} */,
  {32'h41c93e6c, 32'hc3210d70} /* (1, 12, 3) {real, imag} */,
  {32'hc42fd606, 32'hc2beda28} /* (1, 12, 2) {real, imag} */,
  {32'h44a5c934, 32'h4381e1f3} /* (1, 12, 1) {real, imag} */,
  {32'h44563a52, 32'h00000000} /* (1, 12, 0) {real, imag} */,
  {32'h44526876, 32'hc34cab0f} /* (1, 11, 31) {real, imag} */,
  {32'hc3f58278, 32'h4317e0cc} /* (1, 11, 30) {real, imag} */,
  {32'hc264f7a2, 32'hc213a4ca} /* (1, 11, 29) {real, imag} */,
  {32'h42bf4186, 32'hc33bda64} /* (1, 11, 28) {real, imag} */,
  {32'hc23f5f78, 32'h41620f04} /* (1, 11, 27) {real, imag} */,
  {32'h409d2190, 32'h426ae0a8} /* (1, 11, 26) {real, imag} */,
  {32'h429cdc5c, 32'h42216b2a} /* (1, 11, 25) {real, imag} */,
  {32'hc2014e7f, 32'hc202db71} /* (1, 11, 24) {real, imag} */,
  {32'hc29120f6, 32'hc246dc38} /* (1, 11, 23) {real, imag} */,
  {32'h4131b2f2, 32'h421a1eaa} /* (1, 11, 22) {real, imag} */,
  {32'hc2813586, 32'h42479326} /* (1, 11, 21) {real, imag} */,
  {32'h42db3f2e, 32'hc258e401} /* (1, 11, 20) {real, imag} */,
  {32'hc2b01b75, 32'h4188c344} /* (1, 11, 19) {real, imag} */,
  {32'h4168258b, 32'hc001b690} /* (1, 11, 18) {real, imag} */,
  {32'h4142f1fe, 32'hc20903fc} /* (1, 11, 17) {real, imag} */,
  {32'hc16d10b4, 32'h00000000} /* (1, 11, 16) {real, imag} */,
  {32'h4142f1fe, 32'h420903fc} /* (1, 11, 15) {real, imag} */,
  {32'h4168258b, 32'h4001b690} /* (1, 11, 14) {real, imag} */,
  {32'hc2b01b75, 32'hc188c344} /* (1, 11, 13) {real, imag} */,
  {32'h42db3f2e, 32'h4258e401} /* (1, 11, 12) {real, imag} */,
  {32'hc2813586, 32'hc2479326} /* (1, 11, 11) {real, imag} */,
  {32'h4131b2f2, 32'hc21a1eaa} /* (1, 11, 10) {real, imag} */,
  {32'hc29120f6, 32'h4246dc38} /* (1, 11, 9) {real, imag} */,
  {32'hc2014e7f, 32'h4202db71} /* (1, 11, 8) {real, imag} */,
  {32'h429cdc5c, 32'hc2216b2a} /* (1, 11, 7) {real, imag} */,
  {32'h409d2190, 32'hc26ae0a8} /* (1, 11, 6) {real, imag} */,
  {32'hc23f5f78, 32'hc1620f04} /* (1, 11, 5) {real, imag} */,
  {32'h42bf4186, 32'h433bda64} /* (1, 11, 4) {real, imag} */,
  {32'hc264f7a2, 32'h4213a4ca} /* (1, 11, 3) {real, imag} */,
  {32'hc3f58278, 32'hc317e0cc} /* (1, 11, 2) {real, imag} */,
  {32'h44526876, 32'h434cab0f} /* (1, 11, 1) {real, imag} */,
  {32'h43c2300f, 32'h00000000} /* (1, 11, 0) {real, imag} */,
  {32'hc1f3d020, 32'h3f2a6100} /* (1, 10, 31) {real, imag} */,
  {32'h420a342c, 32'h42975d78} /* (1, 10, 30) {real, imag} */,
  {32'hc089a090, 32'hc2a2b410} /* (1, 10, 29) {real, imag} */,
  {32'hc282f9f0, 32'hc2e49640} /* (1, 10, 28) {real, imag} */,
  {32'h4264e923, 32'hc310281a} /* (1, 10, 27) {real, imag} */,
  {32'hc2ba7035, 32'hc0367e1c} /* (1, 10, 26) {real, imag} */,
  {32'h41c7a4a4, 32'h426e9953} /* (1, 10, 25) {real, imag} */,
  {32'h421aa68e, 32'hc11388e3} /* (1, 10, 24) {real, imag} */,
  {32'h41426492, 32'hc197db71} /* (1, 10, 23) {real, imag} */,
  {32'h42cea7e7, 32'h41fbba4e} /* (1, 10, 22) {real, imag} */,
  {32'hc25ea1a9, 32'hc24cc57a} /* (1, 10, 21) {real, imag} */,
  {32'h423120c4, 32'hc1c9a298} /* (1, 10, 20) {real, imag} */,
  {32'hc21cd692, 32'h42a873f2} /* (1, 10, 19) {real, imag} */,
  {32'hc1a2d78c, 32'hc12fcea8} /* (1, 10, 18) {real, imag} */,
  {32'hc209db58, 32'hc12fd1ad} /* (1, 10, 17) {real, imag} */,
  {32'h428424bc, 32'h00000000} /* (1, 10, 16) {real, imag} */,
  {32'hc209db58, 32'h412fd1ad} /* (1, 10, 15) {real, imag} */,
  {32'hc1a2d78c, 32'h412fcea8} /* (1, 10, 14) {real, imag} */,
  {32'hc21cd692, 32'hc2a873f2} /* (1, 10, 13) {real, imag} */,
  {32'h423120c4, 32'h41c9a298} /* (1, 10, 12) {real, imag} */,
  {32'hc25ea1a9, 32'h424cc57a} /* (1, 10, 11) {real, imag} */,
  {32'h42cea7e7, 32'hc1fbba4e} /* (1, 10, 10) {real, imag} */,
  {32'h41426492, 32'h4197db71} /* (1, 10, 9) {real, imag} */,
  {32'h421aa68e, 32'h411388e3} /* (1, 10, 8) {real, imag} */,
  {32'h41c7a4a4, 32'hc26e9953} /* (1, 10, 7) {real, imag} */,
  {32'hc2ba7035, 32'h40367e1c} /* (1, 10, 6) {real, imag} */,
  {32'h4264e923, 32'h4310281a} /* (1, 10, 5) {real, imag} */,
  {32'hc282f9f0, 32'h42e49640} /* (1, 10, 4) {real, imag} */,
  {32'hc089a090, 32'h42a2b410} /* (1, 10, 3) {real, imag} */,
  {32'h420a342c, 32'hc2975d78} /* (1, 10, 2) {real, imag} */,
  {32'hc1f3d020, 32'hbf2a6100} /* (1, 10, 1) {real, imag} */,
  {32'hc35e3766, 32'h00000000} /* (1, 10, 0) {real, imag} */,
  {32'hc43d90c2, 32'h43421f38} /* (1, 9, 31) {real, imag} */,
  {32'h43c23948, 32'hc307a6bc} /* (1, 9, 30) {real, imag} */,
  {32'hc2178059, 32'hc2c63b24} /* (1, 9, 29) {real, imag} */,
  {32'hc3222b1e, 32'hc20c3c6e} /* (1, 9, 28) {real, imag} */,
  {32'h43193dd6, 32'hc2d7bbe9} /* (1, 9, 27) {real, imag} */,
  {32'h416be4c2, 32'hc238cc5f} /* (1, 9, 26) {real, imag} */,
  {32'hc0ddf3ae, 32'h43213d54} /* (1, 9, 25) {real, imag} */,
  {32'h42ce8a86, 32'hc31310ec} /* (1, 9, 24) {real, imag} */,
  {32'h4237e68a, 32'h42c84a50} /* (1, 9, 23) {real, imag} */,
  {32'h421ce4d6, 32'hc1d89f9a} /* (1, 9, 22) {real, imag} */,
  {32'h4273f2df, 32'h410f44e0} /* (1, 9, 21) {real, imag} */,
  {32'hc0d53020, 32'h42d16d9c} /* (1, 9, 20) {real, imag} */,
  {32'h3fb74154, 32'h4044093c} /* (1, 9, 19) {real, imag} */,
  {32'hc2ec723d, 32'hc26ca635} /* (1, 9, 18) {real, imag} */,
  {32'h3fec6640, 32'hc2509f06} /* (1, 9, 17) {real, imag} */,
  {32'hc1ed7306, 32'h00000000} /* (1, 9, 16) {real, imag} */,
  {32'h3fec6640, 32'h42509f06} /* (1, 9, 15) {real, imag} */,
  {32'hc2ec723d, 32'h426ca635} /* (1, 9, 14) {real, imag} */,
  {32'h3fb74154, 32'hc044093c} /* (1, 9, 13) {real, imag} */,
  {32'hc0d53020, 32'hc2d16d9c} /* (1, 9, 12) {real, imag} */,
  {32'h4273f2df, 32'hc10f44e0} /* (1, 9, 11) {real, imag} */,
  {32'h421ce4d6, 32'h41d89f9a} /* (1, 9, 10) {real, imag} */,
  {32'h4237e68a, 32'hc2c84a50} /* (1, 9, 9) {real, imag} */,
  {32'h42ce8a86, 32'h431310ec} /* (1, 9, 8) {real, imag} */,
  {32'hc0ddf3ae, 32'hc3213d54} /* (1, 9, 7) {real, imag} */,
  {32'h416be4c2, 32'h4238cc5f} /* (1, 9, 6) {real, imag} */,
  {32'h43193dd6, 32'h42d7bbe9} /* (1, 9, 5) {real, imag} */,
  {32'hc3222b1e, 32'h420c3c6e} /* (1, 9, 4) {real, imag} */,
  {32'hc2178059, 32'h42c63b24} /* (1, 9, 3) {real, imag} */,
  {32'h43c23948, 32'h4307a6bc} /* (1, 9, 2) {real, imag} */,
  {32'hc43d90c2, 32'hc3421f38} /* (1, 9, 1) {real, imag} */,
  {32'hc43f94c9, 32'h00000000} /* (1, 9, 0) {real, imag} */,
  {32'hc4732e91, 32'h438c30ac} /* (1, 8, 31) {real, imag} */,
  {32'h440dc88c, 32'hc3328475} /* (1, 8, 30) {real, imag} */,
  {32'hc2ae6bcb, 32'hc31aed1e} /* (1, 8, 29) {real, imag} */,
  {32'hc2e1ec15, 32'hc2062be6} /* (1, 8, 28) {real, imag} */,
  {32'h43432e04, 32'h414d1f48} /* (1, 8, 27) {real, imag} */,
  {32'h4283c030, 32'hc257185e} /* (1, 8, 26) {real, imag} */,
  {32'hc23b83ae, 32'hc1852fb0} /* (1, 8, 25) {real, imag} */,
  {32'h42c6359f, 32'hc29b7096} /* (1, 8, 24) {real, imag} */,
  {32'hc13bad50, 32'hbfb5bcc0} /* (1, 8, 23) {real, imag} */,
  {32'h420e51b5, 32'h420ae782} /* (1, 8, 22) {real, imag} */,
  {32'h42e36eee, 32'hc2830649} /* (1, 8, 21) {real, imag} */,
  {32'h42670225, 32'h43191361} /* (1, 8, 20) {real, imag} */,
  {32'hc26b4fb4, 32'h4274a8cc} /* (1, 8, 19) {real, imag} */,
  {32'h4188330a, 32'h42665630} /* (1, 8, 18) {real, imag} */,
  {32'h41b1fa86, 32'h41b8b896} /* (1, 8, 17) {real, imag} */,
  {32'hc1b14df4, 32'h00000000} /* (1, 8, 16) {real, imag} */,
  {32'h41b1fa86, 32'hc1b8b896} /* (1, 8, 15) {real, imag} */,
  {32'h4188330a, 32'hc2665630} /* (1, 8, 14) {real, imag} */,
  {32'hc26b4fb4, 32'hc274a8cc} /* (1, 8, 13) {real, imag} */,
  {32'h42670225, 32'hc3191361} /* (1, 8, 12) {real, imag} */,
  {32'h42e36eee, 32'h42830649} /* (1, 8, 11) {real, imag} */,
  {32'h420e51b5, 32'hc20ae782} /* (1, 8, 10) {real, imag} */,
  {32'hc13bad50, 32'h3fb5bcc0} /* (1, 8, 9) {real, imag} */,
  {32'h42c6359f, 32'h429b7096} /* (1, 8, 8) {real, imag} */,
  {32'hc23b83ae, 32'h41852fb0} /* (1, 8, 7) {real, imag} */,
  {32'h4283c030, 32'h4257185e} /* (1, 8, 6) {real, imag} */,
  {32'h43432e04, 32'hc14d1f48} /* (1, 8, 5) {real, imag} */,
  {32'hc2e1ec15, 32'h42062be6} /* (1, 8, 4) {real, imag} */,
  {32'hc2ae6bcb, 32'h431aed1e} /* (1, 8, 3) {real, imag} */,
  {32'h440dc88c, 32'h43328475} /* (1, 8, 2) {real, imag} */,
  {32'hc4732e91, 32'hc38c30ac} /* (1, 8, 1) {real, imag} */,
  {32'hc45e71ac, 32'h00000000} /* (1, 8, 0) {real, imag} */,
  {32'hc4a3aa57, 32'h43b5fff0} /* (1, 7, 31) {real, imag} */,
  {32'h44344bf3, 32'hc2fb8e7b} /* (1, 7, 30) {real, imag} */,
  {32'h4099c4be, 32'hc317e2b4} /* (1, 7, 29) {real, imag} */,
  {32'hc26ec4fa, 32'hc32c32e6} /* (1, 7, 28) {real, imag} */,
  {32'h43306f01, 32'h42880928} /* (1, 7, 27) {real, imag} */,
  {32'hc16deb08, 32'hc2147e80} /* (1, 7, 26) {real, imag} */,
  {32'hc12b8728, 32'hc1d10fa0} /* (1, 7, 25) {real, imag} */,
  {32'h42fd77b6, 32'hc1c24de0} /* (1, 7, 24) {real, imag} */,
  {32'h425fc218, 32'hc28ca8a7} /* (1, 7, 23) {real, imag} */,
  {32'h420fb492, 32'h41ae4bb1} /* (1, 7, 22) {real, imag} */,
  {32'h431ca136, 32'h41c9faf8} /* (1, 7, 21) {real, imag} */,
  {32'h4278155f, 32'hc19e9dca} /* (1, 7, 20) {real, imag} */,
  {32'h424c0e5a, 32'h422dc515} /* (1, 7, 19) {real, imag} */,
  {32'hc1861f63, 32'h424ad1d9} /* (1, 7, 18) {real, imag} */,
  {32'hc2383f4e, 32'hbfbe9958} /* (1, 7, 17) {real, imag} */,
  {32'hc22b767e, 32'h00000000} /* (1, 7, 16) {real, imag} */,
  {32'hc2383f4e, 32'h3fbe9958} /* (1, 7, 15) {real, imag} */,
  {32'hc1861f63, 32'hc24ad1d9} /* (1, 7, 14) {real, imag} */,
  {32'h424c0e5a, 32'hc22dc515} /* (1, 7, 13) {real, imag} */,
  {32'h4278155f, 32'h419e9dca} /* (1, 7, 12) {real, imag} */,
  {32'h431ca136, 32'hc1c9faf8} /* (1, 7, 11) {real, imag} */,
  {32'h420fb492, 32'hc1ae4bb1} /* (1, 7, 10) {real, imag} */,
  {32'h425fc218, 32'h428ca8a7} /* (1, 7, 9) {real, imag} */,
  {32'h42fd77b6, 32'h41c24de0} /* (1, 7, 8) {real, imag} */,
  {32'hc12b8728, 32'h41d10fa0} /* (1, 7, 7) {real, imag} */,
  {32'hc16deb08, 32'h42147e80} /* (1, 7, 6) {real, imag} */,
  {32'h43306f01, 32'hc2880928} /* (1, 7, 5) {real, imag} */,
  {32'hc26ec4fa, 32'h432c32e6} /* (1, 7, 4) {real, imag} */,
  {32'h4099c4be, 32'h4317e2b4} /* (1, 7, 3) {real, imag} */,
  {32'h44344bf3, 32'h42fb8e7b} /* (1, 7, 2) {real, imag} */,
  {32'hc4a3aa57, 32'hc3b5fff0} /* (1, 7, 1) {real, imag} */,
  {32'hc486b938, 32'h00000000} /* (1, 7, 0) {real, imag} */,
  {32'hc4906a42, 32'h440bb469} /* (1, 6, 31) {real, imag} */,
  {32'h442b783b, 32'hc2e67bf6} /* (1, 6, 30) {real, imag} */,
  {32'h42b9ff45, 32'h3f4a67c0} /* (1, 6, 29) {real, imag} */,
  {32'hc2e70981, 32'hc31917eb} /* (1, 6, 28) {real, imag} */,
  {32'h430bbce8, 32'hc12b56d4} /* (1, 6, 27) {real, imag} */,
  {32'h411ff058, 32'h429455e5} /* (1, 6, 26) {real, imag} */,
  {32'hc263756b, 32'h42f7bcb2} /* (1, 6, 25) {real, imag} */,
  {32'h42dd333d, 32'hc31f7e5f} /* (1, 6, 24) {real, imag} */,
  {32'hc30b600e, 32'hc2200c0c} /* (1, 6, 23) {real, imag} */,
  {32'h40d7d9e8, 32'h430c2074} /* (1, 6, 22) {real, imag} */,
  {32'hc2074a1e, 32'hc248dfb4} /* (1, 6, 21) {real, imag} */,
  {32'hc2b45165, 32'hc052fbb8} /* (1, 6, 20) {real, imag} */,
  {32'h43051c58, 32'h4286c13e} /* (1, 6, 19) {real, imag} */,
  {32'hc25fc3ee, 32'hc2bcc82a} /* (1, 6, 18) {real, imag} */,
  {32'hc241d39e, 32'hc152a80a} /* (1, 6, 17) {real, imag} */,
  {32'h42c13ec3, 32'h00000000} /* (1, 6, 16) {real, imag} */,
  {32'hc241d39e, 32'h4152a80a} /* (1, 6, 15) {real, imag} */,
  {32'hc25fc3ee, 32'h42bcc82a} /* (1, 6, 14) {real, imag} */,
  {32'h43051c58, 32'hc286c13e} /* (1, 6, 13) {real, imag} */,
  {32'hc2b45165, 32'h4052fbb8} /* (1, 6, 12) {real, imag} */,
  {32'hc2074a1e, 32'h4248dfb4} /* (1, 6, 11) {real, imag} */,
  {32'h40d7d9e8, 32'hc30c2074} /* (1, 6, 10) {real, imag} */,
  {32'hc30b600e, 32'h42200c0c} /* (1, 6, 9) {real, imag} */,
  {32'h42dd333d, 32'h431f7e5f} /* (1, 6, 8) {real, imag} */,
  {32'hc263756b, 32'hc2f7bcb2} /* (1, 6, 7) {real, imag} */,
  {32'h411ff058, 32'hc29455e5} /* (1, 6, 6) {real, imag} */,
  {32'h430bbce8, 32'h412b56d4} /* (1, 6, 5) {real, imag} */,
  {32'hc2e70981, 32'h431917eb} /* (1, 6, 4) {real, imag} */,
  {32'h42b9ff45, 32'hbf4a67c0} /* (1, 6, 3) {real, imag} */,
  {32'h442b783b, 32'h42e67bf6} /* (1, 6, 2) {real, imag} */,
  {32'hc4906a42, 32'hc40bb469} /* (1, 6, 1) {real, imag} */,
  {32'hc47ce040, 32'h00000000} /* (1, 6, 0) {real, imag} */,
  {32'hc460b8f4, 32'h447e147b} /* (1, 5, 31) {real, imag} */,
  {32'h42d5c1c0, 32'hc35c8d72} /* (1, 5, 30) {real, imag} */,
  {32'h433c1752, 32'hc1ad8f5b} /* (1, 5, 29) {real, imag} */,
  {32'hc30aa347, 32'hc1f4eb60} /* (1, 5, 28) {real, imag} */,
  {32'h433f2a7a, 32'hc22c07e7} /* (1, 5, 27) {real, imag} */,
  {32'hc0f57820, 32'hc0ad5f00} /* (1, 5, 26) {real, imag} */,
  {32'hc0b7a578, 32'h42f47826} /* (1, 5, 25) {real, imag} */,
  {32'h432c48d4, 32'hc2652ff5} /* (1, 5, 24) {real, imag} */,
  {32'hc240aaac, 32'hc27d6e89} /* (1, 5, 23) {real, imag} */,
  {32'hc20ba544, 32'hc1f908d7} /* (1, 5, 22) {real, imag} */,
  {32'h41ef9650, 32'h41c7fa57} /* (1, 5, 21) {real, imag} */,
  {32'h42116a47, 32'h41e8781a} /* (1, 5, 20) {real, imag} */,
  {32'h427026d0, 32'h41a87a42} /* (1, 5, 19) {real, imag} */,
  {32'h425d5842, 32'hc2bbd289} /* (1, 5, 18) {real, imag} */,
  {32'hc23cc4a6, 32'h41f26377} /* (1, 5, 17) {real, imag} */,
  {32'hc280deb2, 32'h00000000} /* (1, 5, 16) {real, imag} */,
  {32'hc23cc4a6, 32'hc1f26377} /* (1, 5, 15) {real, imag} */,
  {32'h425d5842, 32'h42bbd289} /* (1, 5, 14) {real, imag} */,
  {32'h427026d0, 32'hc1a87a42} /* (1, 5, 13) {real, imag} */,
  {32'h42116a47, 32'hc1e8781a} /* (1, 5, 12) {real, imag} */,
  {32'h41ef9650, 32'hc1c7fa57} /* (1, 5, 11) {real, imag} */,
  {32'hc20ba544, 32'h41f908d7} /* (1, 5, 10) {real, imag} */,
  {32'hc240aaac, 32'h427d6e89} /* (1, 5, 9) {real, imag} */,
  {32'h432c48d4, 32'h42652ff5} /* (1, 5, 8) {real, imag} */,
  {32'hc0b7a578, 32'hc2f47826} /* (1, 5, 7) {real, imag} */,
  {32'hc0f57820, 32'h40ad5f00} /* (1, 5, 6) {real, imag} */,
  {32'h433f2a7a, 32'h422c07e7} /* (1, 5, 5) {real, imag} */,
  {32'hc30aa347, 32'h41f4eb60} /* (1, 5, 4) {real, imag} */,
  {32'h433c1752, 32'h41ad8f5b} /* (1, 5, 3) {real, imag} */,
  {32'h42d5c1c0, 32'h435c8d72} /* (1, 5, 2) {real, imag} */,
  {32'hc460b8f4, 32'hc47e147b} /* (1, 5, 1) {real, imag} */,
  {32'hc495a8fc, 32'h00000000} /* (1, 5, 0) {real, imag} */,
  {32'hc4462304, 32'h44a25e3c} /* (1, 4, 31) {real, imag} */,
  {32'hc3896f0c, 32'hc38c3bc5} /* (1, 4, 30) {real, imag} */,
  {32'h435f5c22, 32'hc30f3ec1} /* (1, 4, 29) {real, imag} */,
  {32'h3fc96780, 32'hc36e66c3} /* (1, 4, 28) {real, imag} */,
  {32'h42a9a29a, 32'h41c5fc44} /* (1, 4, 27) {real, imag} */,
  {32'h422e4f31, 32'hc00a9d50} /* (1, 4, 26) {real, imag} */,
  {32'h42a8ee32, 32'hc1125978} /* (1, 4, 25) {real, imag} */,
  {32'hc24b99c9, 32'hc184b836} /* (1, 4, 24) {real, imag} */,
  {32'h42b534b2, 32'h40988c5c} /* (1, 4, 23) {real, imag} */,
  {32'hc14a8dee, 32'hc27dc711} /* (1, 4, 22) {real, imag} */,
  {32'h42731bc1, 32'h42877d07} /* (1, 4, 21) {real, imag} */,
  {32'h40582142, 32'hc20290ab} /* (1, 4, 20) {real, imag} */,
  {32'hc212b90a, 32'hc20f7ba6} /* (1, 4, 19) {real, imag} */,
  {32'h42890c95, 32'h4183277f} /* (1, 4, 18) {real, imag} */,
  {32'h4206458d, 32'h41dc0fff} /* (1, 4, 17) {real, imag} */,
  {32'h41e35905, 32'h00000000} /* (1, 4, 16) {real, imag} */,
  {32'h4206458d, 32'hc1dc0fff} /* (1, 4, 15) {real, imag} */,
  {32'h42890c95, 32'hc183277f} /* (1, 4, 14) {real, imag} */,
  {32'hc212b90a, 32'h420f7ba6} /* (1, 4, 13) {real, imag} */,
  {32'h40582142, 32'h420290ab} /* (1, 4, 12) {real, imag} */,
  {32'h42731bc1, 32'hc2877d07} /* (1, 4, 11) {real, imag} */,
  {32'hc14a8dee, 32'h427dc711} /* (1, 4, 10) {real, imag} */,
  {32'h42b534b2, 32'hc0988c5c} /* (1, 4, 9) {real, imag} */,
  {32'hc24b99c9, 32'h4184b836} /* (1, 4, 8) {real, imag} */,
  {32'h42a8ee32, 32'h41125978} /* (1, 4, 7) {real, imag} */,
  {32'h422e4f31, 32'h400a9d50} /* (1, 4, 6) {real, imag} */,
  {32'h42a9a29a, 32'hc1c5fc44} /* (1, 4, 5) {real, imag} */,
  {32'h3fc96780, 32'h436e66c3} /* (1, 4, 4) {real, imag} */,
  {32'h435f5c22, 32'h430f3ec1} /* (1, 4, 3) {real, imag} */,
  {32'hc3896f0c, 32'h438c3bc5} /* (1, 4, 2) {real, imag} */,
  {32'hc4462304, 32'hc4a25e3c} /* (1, 4, 1) {real, imag} */,
  {32'hc49f4694, 32'h00000000} /* (1, 4, 0) {real, imag} */,
  {32'hc42af1c2, 32'h44b1a81e} /* (1, 3, 31) {real, imag} */,
  {32'hc381fe95, 32'hc3ff2a62} /* (1, 3, 30) {real, imag} */,
  {32'h438563eb, 32'h40559710} /* (1, 3, 29) {real, imag} */,
  {32'h425f15e6, 32'hc3254ecf} /* (1, 3, 28) {real, imag} */,
  {32'h4256d51a, 32'h43295118} /* (1, 3, 27) {real, imag} */,
  {32'h42d57b12, 32'hc23cc858} /* (1, 3, 26) {real, imag} */,
  {32'hc23c365c, 32'h414537fc} /* (1, 3, 25) {real, imag} */,
  {32'hc1c7c8a8, 32'h41ea140e} /* (1, 3, 24) {real, imag} */,
  {32'h42b1407c, 32'hc2865de2} /* (1, 3, 23) {real, imag} */,
  {32'h4266cc1e, 32'h4281ab5f} /* (1, 3, 22) {real, imag} */,
  {32'hc290de06, 32'h41a3dfb4} /* (1, 3, 21) {real, imag} */,
  {32'hc2e664a0, 32'h4105500c} /* (1, 3, 20) {real, imag} */,
  {32'hc0961ce0, 32'h418b91f2} /* (1, 3, 19) {real, imag} */,
  {32'hc1ff5bf8, 32'hc2435aee} /* (1, 3, 18) {real, imag} */,
  {32'h415b1c83, 32'hc194abd8} /* (1, 3, 17) {real, imag} */,
  {32'h427e5f7d, 32'h00000000} /* (1, 3, 16) {real, imag} */,
  {32'h415b1c83, 32'h4194abd8} /* (1, 3, 15) {real, imag} */,
  {32'hc1ff5bf8, 32'h42435aee} /* (1, 3, 14) {real, imag} */,
  {32'hc0961ce0, 32'hc18b91f2} /* (1, 3, 13) {real, imag} */,
  {32'hc2e664a0, 32'hc105500c} /* (1, 3, 12) {real, imag} */,
  {32'hc290de06, 32'hc1a3dfb4} /* (1, 3, 11) {real, imag} */,
  {32'h4266cc1e, 32'hc281ab5f} /* (1, 3, 10) {real, imag} */,
  {32'h42b1407c, 32'h42865de2} /* (1, 3, 9) {real, imag} */,
  {32'hc1c7c8a8, 32'hc1ea140e} /* (1, 3, 8) {real, imag} */,
  {32'hc23c365c, 32'hc14537fc} /* (1, 3, 7) {real, imag} */,
  {32'h42d57b12, 32'h423cc858} /* (1, 3, 6) {real, imag} */,
  {32'h4256d51a, 32'hc3295118} /* (1, 3, 5) {real, imag} */,
  {32'h425f15e6, 32'h43254ecf} /* (1, 3, 4) {real, imag} */,
  {32'h438563eb, 32'hc0559710} /* (1, 3, 3) {real, imag} */,
  {32'hc381fe95, 32'h43ff2a62} /* (1, 3, 2) {real, imag} */,
  {32'hc42af1c2, 32'hc4b1a81e} /* (1, 3, 1) {real, imag} */,
  {32'hc490a92e, 32'h00000000} /* (1, 3, 0) {real, imag} */,
  {32'hc465c8b5, 32'h44a92c60} /* (1, 2, 31) {real, imag} */,
  {32'hc3ebb10a, 32'hc40fb3a0} /* (1, 2, 30) {real, imag} */,
  {32'h4381f710, 32'h4212f3ef} /* (1, 2, 29) {real, imag} */,
  {32'h400e2ba0, 32'hc380db88} /* (1, 2, 28) {real, imag} */,
  {32'h4334d18c, 32'h42b631f6} /* (1, 2, 27) {real, imag} */,
  {32'h40257a10, 32'hc24680fe} /* (1, 2, 26) {real, imag} */,
  {32'hc204fc1f, 32'h419a7bae} /* (1, 2, 25) {real, imag} */,
  {32'hc2cf7467, 32'h3ee47f80} /* (1, 2, 24) {real, imag} */,
  {32'hc3219510, 32'hc307a5d8} /* (1, 2, 23) {real, imag} */,
  {32'h42abd29e, 32'hc24d394e} /* (1, 2, 22) {real, imag} */,
  {32'h42c93eac, 32'hc1224534} /* (1, 2, 21) {real, imag} */,
  {32'h42e1eb50, 32'hc291069a} /* (1, 2, 20) {real, imag} */,
  {32'hc16215e6, 32'h404f385c} /* (1, 2, 19) {real, imag} */,
  {32'hc295a670, 32'hc2ee53c9} /* (1, 2, 18) {real, imag} */,
  {32'h41f1354c, 32'hc1b61fea} /* (1, 2, 17) {real, imag} */,
  {32'hc11d5804, 32'h00000000} /* (1, 2, 16) {real, imag} */,
  {32'h41f1354c, 32'h41b61fea} /* (1, 2, 15) {real, imag} */,
  {32'hc295a670, 32'h42ee53c9} /* (1, 2, 14) {real, imag} */,
  {32'hc16215e6, 32'hc04f385c} /* (1, 2, 13) {real, imag} */,
  {32'h42e1eb50, 32'h4291069a} /* (1, 2, 12) {real, imag} */,
  {32'h42c93eac, 32'h41224534} /* (1, 2, 11) {real, imag} */,
  {32'h42abd29e, 32'h424d394e} /* (1, 2, 10) {real, imag} */,
  {32'hc3219510, 32'h4307a5d8} /* (1, 2, 9) {real, imag} */,
  {32'hc2cf7467, 32'hbee47f80} /* (1, 2, 8) {real, imag} */,
  {32'hc204fc1f, 32'hc19a7bae} /* (1, 2, 7) {real, imag} */,
  {32'h40257a10, 32'h424680fe} /* (1, 2, 6) {real, imag} */,
  {32'h4334d18c, 32'hc2b631f6} /* (1, 2, 5) {real, imag} */,
  {32'h400e2ba0, 32'h4380db88} /* (1, 2, 4) {real, imag} */,
  {32'h4381f710, 32'hc212f3ef} /* (1, 2, 3) {real, imag} */,
  {32'hc3ebb10a, 32'h440fb3a0} /* (1, 2, 2) {real, imag} */,
  {32'hc465c8b5, 32'hc4a92c60} /* (1, 2, 1) {real, imag} */,
  {32'hc46e94e9, 32'h00000000} /* (1, 2, 0) {real, imag} */,
  {32'hc45a7438, 32'h448d5d3a} /* (1, 1, 31) {real, imag} */,
  {32'hc3aaea9c, 32'hc4236a54} /* (1, 1, 30) {real, imag} */,
  {32'h436eb8da, 32'hc1f57be9} /* (1, 1, 29) {real, imag} */,
  {32'h4201b0ca, 32'hc372e8ce} /* (1, 1, 28) {real, imag} */,
  {32'h438628cc, 32'h4342b51a} /* (1, 1, 27) {real, imag} */,
  {32'h4206682e, 32'h42c483f8} /* (1, 1, 26) {real, imag} */,
  {32'hc2866f60, 32'h41fbf318} /* (1, 1, 25) {real, imag} */,
  {32'hc2806a02, 32'h41e2573a} /* (1, 1, 24) {real, imag} */,
  {32'hc26815f2, 32'hc2cc8220} /* (1, 1, 23) {real, imag} */,
  {32'h400ae480, 32'hc2725a9b} /* (1, 1, 22) {real, imag} */,
  {32'h413a61d4, 32'hc288e3fb} /* (1, 1, 21) {real, imag} */,
  {32'h42aadc4d, 32'h41b69f19} /* (1, 1, 20) {real, imag} */,
  {32'h41638184, 32'h4084d8b0} /* (1, 1, 19) {real, imag} */,
  {32'hc0f68a82, 32'h3ff251d0} /* (1, 1, 18) {real, imag} */,
  {32'h3f8168e0, 32'h421e676e} /* (1, 1, 17) {real, imag} */,
  {32'hc2cafe9e, 32'h00000000} /* (1, 1, 16) {real, imag} */,
  {32'h3f8168e0, 32'hc21e676e} /* (1, 1, 15) {real, imag} */,
  {32'hc0f68a82, 32'hbff251d0} /* (1, 1, 14) {real, imag} */,
  {32'h41638184, 32'hc084d8b0} /* (1, 1, 13) {real, imag} */,
  {32'h42aadc4d, 32'hc1b69f19} /* (1, 1, 12) {real, imag} */,
  {32'h413a61d4, 32'h4288e3fb} /* (1, 1, 11) {real, imag} */,
  {32'h400ae480, 32'h42725a9b} /* (1, 1, 10) {real, imag} */,
  {32'hc26815f2, 32'h42cc8220} /* (1, 1, 9) {real, imag} */,
  {32'hc2806a02, 32'hc1e2573a} /* (1, 1, 8) {real, imag} */,
  {32'hc2866f60, 32'hc1fbf318} /* (1, 1, 7) {real, imag} */,
  {32'h4206682e, 32'hc2c483f8} /* (1, 1, 6) {real, imag} */,
  {32'h438628cc, 32'hc342b51a} /* (1, 1, 5) {real, imag} */,
  {32'h4201b0ca, 32'h4372e8ce} /* (1, 1, 4) {real, imag} */,
  {32'h436eb8da, 32'h41f57be9} /* (1, 1, 3) {real, imag} */,
  {32'hc3aaea9c, 32'h44236a54} /* (1, 1, 2) {real, imag} */,
  {32'hc45a7438, 32'hc48d5d3a} /* (1, 1, 1) {real, imag} */,
  {32'hc41b44da, 32'h00000000} /* (1, 1, 0) {real, imag} */,
  {32'hc439d1e3, 32'h443c5560} /* (1, 0, 31) {real, imag} */,
  {32'hc2ea4aa0, 32'hc3d59685} /* (1, 0, 30) {real, imag} */,
  {32'h425e0f24, 32'hc25b6ffc} /* (1, 0, 29) {real, imag} */,
  {32'h3f07f300, 32'hc2cb3860} /* (1, 0, 28) {real, imag} */,
  {32'h42e6bf5a, 32'h422a7042} /* (1, 0, 27) {real, imag} */,
  {32'h41207f60, 32'hc25eaa06} /* (1, 0, 26) {real, imag} */,
  {32'hc28d7372, 32'h42758db3} /* (1, 0, 25) {real, imag} */,
  {32'h41a1a23e, 32'h4257197c} /* (1, 0, 24) {real, imag} */,
  {32'h42e50854, 32'hc2ee28ce} /* (1, 0, 23) {real, imag} */,
  {32'hc22fad34, 32'h427f15ff} /* (1, 0, 22) {real, imag} */,
  {32'hc23755c6, 32'h42564520} /* (1, 0, 21) {real, imag} */,
  {32'h4020b670, 32'h41de09fd} /* (1, 0, 20) {real, imag} */,
  {32'h41124aa8, 32'hc2729dd9} /* (1, 0, 19) {real, imag} */,
  {32'hc1aaabd4, 32'h3fccd848} /* (1, 0, 18) {real, imag} */,
  {32'h41977076, 32'h413518e1} /* (1, 0, 17) {real, imag} */,
  {32'h418ca216, 32'h00000000} /* (1, 0, 16) {real, imag} */,
  {32'h41977076, 32'hc13518e1} /* (1, 0, 15) {real, imag} */,
  {32'hc1aaabd4, 32'hbfccd848} /* (1, 0, 14) {real, imag} */,
  {32'h41124aa8, 32'h42729dd9} /* (1, 0, 13) {real, imag} */,
  {32'h4020b670, 32'hc1de09fd} /* (1, 0, 12) {real, imag} */,
  {32'hc23755c6, 32'hc2564520} /* (1, 0, 11) {real, imag} */,
  {32'hc22fad34, 32'hc27f15ff} /* (1, 0, 10) {real, imag} */,
  {32'h42e50854, 32'h42ee28ce} /* (1, 0, 9) {real, imag} */,
  {32'h41a1a23e, 32'hc257197c} /* (1, 0, 8) {real, imag} */,
  {32'hc28d7372, 32'hc2758db3} /* (1, 0, 7) {real, imag} */,
  {32'h41207f60, 32'h425eaa06} /* (1, 0, 6) {real, imag} */,
  {32'h42e6bf5a, 32'hc22a7042} /* (1, 0, 5) {real, imag} */,
  {32'h3f07f300, 32'h42cb3860} /* (1, 0, 4) {real, imag} */,
  {32'h425e0f24, 32'h425b6ffc} /* (1, 0, 3) {real, imag} */,
  {32'hc2ea4aa0, 32'h43d59685} /* (1, 0, 2) {real, imag} */,
  {32'hc439d1e3, 32'hc43c5560} /* (1, 0, 1) {real, imag} */,
  {32'hc3ec9a39, 32'h00000000} /* (1, 0, 0) {real, imag} */,
  {32'hc3c7693c, 32'h431c1ee2} /* (0, 31, 31) {real, imag} */,
  {32'hc007d080, 32'hc1f251bc} /* (0, 31, 30) {real, imag} */,
  {32'h42ed8fce, 32'h4274e5df} /* (0, 31, 29) {real, imag} */,
  {32'h428a77aa, 32'h41b4377c} /* (0, 31, 28) {real, imag} */,
  {32'h42ed7b1e, 32'hc126e4fa} /* (0, 31, 27) {real, imag} */,
  {32'h4197f6ee, 32'hc29f0477} /* (0, 31, 26) {real, imag} */,
  {32'hc2290855, 32'hc10af7d8} /* (0, 31, 25) {real, imag} */,
  {32'hc2911129, 32'hc2502d4f} /* (0, 31, 24) {real, imag} */,
  {32'hc1e4010a, 32'hc1b7c129} /* (0, 31, 23) {real, imag} */,
  {32'hc241b0d7, 32'h424f5c56} /* (0, 31, 22) {real, imag} */,
  {32'hc0b5c2ac, 32'h41749336} /* (0, 31, 21) {real, imag} */,
  {32'h41d40672, 32'h42458a7c} /* (0, 31, 20) {real, imag} */,
  {32'hc01812e0, 32'hc1ec5e0f} /* (0, 31, 19) {real, imag} */,
  {32'h418e0bf6, 32'hc182e8a4} /* (0, 31, 18) {real, imag} */,
  {32'h40793ce0, 32'hbea3be80} /* (0, 31, 17) {real, imag} */,
  {32'hc1082c30, 32'h00000000} /* (0, 31, 16) {real, imag} */,
  {32'h40793ce0, 32'h3ea3be80} /* (0, 31, 15) {real, imag} */,
  {32'h418e0bf6, 32'h4182e8a4} /* (0, 31, 14) {real, imag} */,
  {32'hc01812e0, 32'h41ec5e0f} /* (0, 31, 13) {real, imag} */,
  {32'h41d40672, 32'hc2458a7c} /* (0, 31, 12) {real, imag} */,
  {32'hc0b5c2ac, 32'hc1749336} /* (0, 31, 11) {real, imag} */,
  {32'hc241b0d7, 32'hc24f5c56} /* (0, 31, 10) {real, imag} */,
  {32'hc1e4010a, 32'h41b7c129} /* (0, 31, 9) {real, imag} */,
  {32'hc2911129, 32'h42502d4f} /* (0, 31, 8) {real, imag} */,
  {32'hc2290855, 32'h410af7d8} /* (0, 31, 7) {real, imag} */,
  {32'h4197f6ee, 32'h429f0477} /* (0, 31, 6) {real, imag} */,
  {32'h42ed7b1e, 32'h4126e4fa} /* (0, 31, 5) {real, imag} */,
  {32'h428a77aa, 32'hc1b4377c} /* (0, 31, 4) {real, imag} */,
  {32'h42ed8fce, 32'hc274e5df} /* (0, 31, 3) {real, imag} */,
  {32'hc007d080, 32'h41f251bc} /* (0, 31, 2) {real, imag} */,
  {32'hc3c7693c, 32'hc31c1ee2} /* (0, 31, 1) {real, imag} */,
  {32'hc39199ed, 32'h00000000} /* (0, 31, 0) {real, imag} */,
  {32'hc401f914, 32'h422fa970} /* (0, 30, 31) {real, imag} */,
  {32'h432d56bd, 32'hc19a74c4} /* (0, 30, 30) {real, imag} */,
  {32'h42cf9ffc, 32'hc1a9842e} /* (0, 30, 29) {real, imag} */,
  {32'h42abca0c, 32'h41f4cf7e} /* (0, 30, 28) {real, imag} */,
  {32'h42ced7b0, 32'h422bce3e} /* (0, 30, 27) {real, imag} */,
  {32'h426c35b3, 32'hc212b3e2} /* (0, 30, 26) {real, imag} */,
  {32'hc285a5ae, 32'h412277d0} /* (0, 30, 25) {real, imag} */,
  {32'hc21433b8, 32'h418238dc} /* (0, 30, 24) {real, imag} */,
  {32'hc224fcf6, 32'h4230fb17} /* (0, 30, 23) {real, imag} */,
  {32'h42762d8c, 32'h4285f620} /* (0, 30, 22) {real, imag} */,
  {32'h41dfd5a3, 32'h41d101f0} /* (0, 30, 21) {real, imag} */,
  {32'h3f966f48, 32'h42dadf9c} /* (0, 30, 20) {real, imag} */,
  {32'hc1bd8169, 32'h414ea566} /* (0, 30, 19) {real, imag} */,
  {32'h420479e1, 32'h40da2e28} /* (0, 30, 18) {real, imag} */,
  {32'h40ce6c30, 32'h416c23f2} /* (0, 30, 17) {real, imag} */,
  {32'h41ad90a7, 32'h00000000} /* (0, 30, 16) {real, imag} */,
  {32'h40ce6c30, 32'hc16c23f2} /* (0, 30, 15) {real, imag} */,
  {32'h420479e1, 32'hc0da2e28} /* (0, 30, 14) {real, imag} */,
  {32'hc1bd8169, 32'hc14ea566} /* (0, 30, 13) {real, imag} */,
  {32'h3f966f48, 32'hc2dadf9c} /* (0, 30, 12) {real, imag} */,
  {32'h41dfd5a3, 32'hc1d101f0} /* (0, 30, 11) {real, imag} */,
  {32'h42762d8c, 32'hc285f620} /* (0, 30, 10) {real, imag} */,
  {32'hc224fcf6, 32'hc230fb17} /* (0, 30, 9) {real, imag} */,
  {32'hc21433b8, 32'hc18238dc} /* (0, 30, 8) {real, imag} */,
  {32'hc285a5ae, 32'hc12277d0} /* (0, 30, 7) {real, imag} */,
  {32'h426c35b3, 32'h4212b3e2} /* (0, 30, 6) {real, imag} */,
  {32'h42ced7b0, 32'hc22bce3e} /* (0, 30, 5) {real, imag} */,
  {32'h42abca0c, 32'hc1f4cf7e} /* (0, 30, 4) {real, imag} */,
  {32'h42cf9ffc, 32'h41a9842e} /* (0, 30, 3) {real, imag} */,
  {32'h432d56bd, 32'h419a74c4} /* (0, 30, 2) {real, imag} */,
  {32'hc401f914, 32'hc22fa970} /* (0, 30, 1) {real, imag} */,
  {32'hc3c59b17, 32'h00000000} /* (0, 30, 0) {real, imag} */,
  {32'hc41fb971, 32'h420cbcc0} /* (0, 29, 31) {real, imag} */,
  {32'h438eccbc, 32'hc225f8b6} /* (0, 29, 30) {real, imag} */,
  {32'h41cc8f7c, 32'h421ecc6e} /* (0, 29, 29) {real, imag} */,
  {32'hc208d5b2, 32'h4221ed47} /* (0, 29, 28) {real, imag} */,
  {32'h426b195e, 32'h3e030c00} /* (0, 29, 27) {real, imag} */,
  {32'h42674c56, 32'h41f79e71} /* (0, 29, 26) {real, imag} */,
  {32'hc2297c0f, 32'hc221bbec} /* (0, 29, 25) {real, imag} */,
  {32'h3df12800, 32'hc1179292} /* (0, 29, 24) {real, imag} */,
  {32'hc010c63c, 32'h41659160} /* (0, 29, 23) {real, imag} */,
  {32'hc1a32771, 32'h42b024e7} /* (0, 29, 22) {real, imag} */,
  {32'hc0ecb038, 32'hc188d813} /* (0, 29, 21) {real, imag} */,
  {32'h41f655fa, 32'h42a8dd5a} /* (0, 29, 20) {real, imag} */,
  {32'hc15769e4, 32'h422b09f4} /* (0, 29, 19) {real, imag} */,
  {32'h419f2260, 32'hc17e1d0a} /* (0, 29, 18) {real, imag} */,
  {32'hc1807490, 32'hbfedd800} /* (0, 29, 17) {real, imag} */,
  {32'h422363c4, 32'h00000000} /* (0, 29, 16) {real, imag} */,
  {32'hc1807490, 32'h3fedd800} /* (0, 29, 15) {real, imag} */,
  {32'h419f2260, 32'h417e1d0a} /* (0, 29, 14) {real, imag} */,
  {32'hc15769e4, 32'hc22b09f4} /* (0, 29, 13) {real, imag} */,
  {32'h41f655fa, 32'hc2a8dd5a} /* (0, 29, 12) {real, imag} */,
  {32'hc0ecb038, 32'h4188d813} /* (0, 29, 11) {real, imag} */,
  {32'hc1a32771, 32'hc2b024e7} /* (0, 29, 10) {real, imag} */,
  {32'hc010c63c, 32'hc1659160} /* (0, 29, 9) {real, imag} */,
  {32'h3df12800, 32'h41179292} /* (0, 29, 8) {real, imag} */,
  {32'hc2297c0f, 32'h4221bbec} /* (0, 29, 7) {real, imag} */,
  {32'h42674c56, 32'hc1f79e71} /* (0, 29, 6) {real, imag} */,
  {32'h426b195e, 32'hbe030c00} /* (0, 29, 5) {real, imag} */,
  {32'hc208d5b2, 32'hc221ed47} /* (0, 29, 4) {real, imag} */,
  {32'h41cc8f7c, 32'hc21ecc6e} /* (0, 29, 3) {real, imag} */,
  {32'h438eccbc, 32'h4225f8b6} /* (0, 29, 2) {real, imag} */,
  {32'hc41fb971, 32'hc20cbcc0} /* (0, 29, 1) {real, imag} */,
  {32'hc3c1ca78, 32'h00000000} /* (0, 29, 0) {real, imag} */,
  {32'hc4325e9e, 32'hc12a2c80} /* (0, 28, 31) {real, imag} */,
  {32'h43519199, 32'h4121866c} /* (0, 28, 30) {real, imag} */,
  {32'h4053b670, 32'h40729570} /* (0, 28, 29) {real, imag} */,
  {32'hc24e88e3, 32'h42faf8d9} /* (0, 28, 28) {real, imag} */,
  {32'h432dd147, 32'hc239116e} /* (0, 28, 27) {real, imag} */,
  {32'h3f896008, 32'h422c43b0} /* (0, 28, 26) {real, imag} */,
  {32'hc1c4acaa, 32'hc116ddcf} /* (0, 28, 25) {real, imag} */,
  {32'h4222fe04, 32'hc2cdda7b} /* (0, 28, 24) {real, imag} */,
  {32'hbff97960, 32'hbfe1cd54} /* (0, 28, 23) {real, imag} */,
  {32'hc1b55427, 32'h4129972d} /* (0, 28, 22) {real, imag} */,
  {32'hc1c86dd0, 32'h4276e3ea} /* (0, 28, 21) {real, imag} */,
  {32'hbf1ef610, 32'h4229b12c} /* (0, 28, 20) {real, imag} */,
  {32'hc19ff3ae, 32'hc248e538} /* (0, 28, 19) {real, imag} */,
  {32'h41248dd8, 32'hc26f3a6d} /* (0, 28, 18) {real, imag} */,
  {32'hc1253012, 32'hc151f96a} /* (0, 28, 17) {real, imag} */,
  {32'h40ab76ae, 32'h00000000} /* (0, 28, 16) {real, imag} */,
  {32'hc1253012, 32'h4151f96a} /* (0, 28, 15) {real, imag} */,
  {32'h41248dd8, 32'h426f3a6d} /* (0, 28, 14) {real, imag} */,
  {32'hc19ff3ae, 32'h4248e538} /* (0, 28, 13) {real, imag} */,
  {32'hbf1ef610, 32'hc229b12c} /* (0, 28, 12) {real, imag} */,
  {32'hc1c86dd0, 32'hc276e3ea} /* (0, 28, 11) {real, imag} */,
  {32'hc1b55427, 32'hc129972d} /* (0, 28, 10) {real, imag} */,
  {32'hbff97960, 32'h3fe1cd54} /* (0, 28, 9) {real, imag} */,
  {32'h4222fe04, 32'h42cdda7b} /* (0, 28, 8) {real, imag} */,
  {32'hc1c4acaa, 32'h4116ddcf} /* (0, 28, 7) {real, imag} */,
  {32'h3f896008, 32'hc22c43b0} /* (0, 28, 6) {real, imag} */,
  {32'h432dd147, 32'h4239116e} /* (0, 28, 5) {real, imag} */,
  {32'hc24e88e3, 32'hc2faf8d9} /* (0, 28, 4) {real, imag} */,
  {32'h4053b670, 32'hc0729570} /* (0, 28, 3) {real, imag} */,
  {32'h43519199, 32'hc121866c} /* (0, 28, 2) {real, imag} */,
  {32'hc4325e9e, 32'h412a2c80} /* (0, 28, 1) {real, imag} */,
  {32'hc3915680, 32'h00000000} /* (0, 28, 0) {real, imag} */,
  {32'hc42b8939, 32'h428acae0} /* (0, 27, 31) {real, imag} */,
  {32'h433a8d1e, 32'h426d0a00} /* (0, 27, 30) {real, imag} */,
  {32'h40ddf218, 32'hc26adaf9} /* (0, 27, 29) {real, imag} */,
  {32'hc1b6bdd2, 32'h430155ba} /* (0, 27, 28) {real, imag} */,
  {32'h42b51949, 32'hc1eb3028} /* (0, 27, 27) {real, imag} */,
  {32'h4110ff94, 32'h4190e5d2} /* (0, 27, 26) {real, imag} */,
  {32'hc2468046, 32'hc18b9926} /* (0, 27, 25) {real, imag} */,
  {32'hc0e8fc76, 32'h40b3a2bc} /* (0, 27, 24) {real, imag} */,
  {32'h417ce8c4, 32'hc2ae8e96} /* (0, 27, 23) {real, imag} */,
  {32'hc24eab14, 32'hc07a0c00} /* (0, 27, 22) {real, imag} */,
  {32'h4250ba80, 32'hc018ef00} /* (0, 27, 21) {real, imag} */,
  {32'hc198ad5a, 32'h400efaa0} /* (0, 27, 20) {real, imag} */,
  {32'h41c31608, 32'hc1c6d1b6} /* (0, 27, 19) {real, imag} */,
  {32'hbfeebd20, 32'hc21c57bd} /* (0, 27, 18) {real, imag} */,
  {32'hc0bf58fe, 32'h420bf8e4} /* (0, 27, 17) {real, imag} */,
  {32'hc2a084a2, 32'h00000000} /* (0, 27, 16) {real, imag} */,
  {32'hc0bf58fe, 32'hc20bf8e4} /* (0, 27, 15) {real, imag} */,
  {32'hbfeebd20, 32'h421c57bd} /* (0, 27, 14) {real, imag} */,
  {32'h41c31608, 32'h41c6d1b6} /* (0, 27, 13) {real, imag} */,
  {32'hc198ad5a, 32'hc00efaa0} /* (0, 27, 12) {real, imag} */,
  {32'h4250ba80, 32'h4018ef00} /* (0, 27, 11) {real, imag} */,
  {32'hc24eab14, 32'h407a0c00} /* (0, 27, 10) {real, imag} */,
  {32'h417ce8c4, 32'h42ae8e96} /* (0, 27, 9) {real, imag} */,
  {32'hc0e8fc76, 32'hc0b3a2bc} /* (0, 27, 8) {real, imag} */,
  {32'hc2468046, 32'h418b9926} /* (0, 27, 7) {real, imag} */,
  {32'h4110ff94, 32'hc190e5d2} /* (0, 27, 6) {real, imag} */,
  {32'h42b51949, 32'h41eb3028} /* (0, 27, 5) {real, imag} */,
  {32'hc1b6bdd2, 32'hc30155ba} /* (0, 27, 4) {real, imag} */,
  {32'h40ddf218, 32'h426adaf9} /* (0, 27, 3) {real, imag} */,
  {32'h433a8d1e, 32'hc26d0a00} /* (0, 27, 2) {real, imag} */,
  {32'hc42b8939, 32'hc28acae0} /* (0, 27, 1) {real, imag} */,
  {32'hc388f38b, 32'h00000000} /* (0, 27, 0) {real, imag} */,
  {32'hc4496816, 32'h427bd300} /* (0, 26, 31) {real, imag} */,
  {32'h433c427b, 32'h42aec14d} /* (0, 26, 30) {real, imag} */,
  {32'hc212b92c, 32'hc229c27f} /* (0, 26, 29) {real, imag} */,
  {32'hc2fa53e6, 32'h42e19571} /* (0, 26, 28) {real, imag} */,
  {32'h4311c5c2, 32'hc20018cf} /* (0, 26, 27) {real, imag} */,
  {32'h41ca84b3, 32'hc0a2f3c0} /* (0, 26, 26) {real, imag} */,
  {32'h41e0f145, 32'h428be12f} /* (0, 26, 25) {real, imag} */,
  {32'h4255470a, 32'hc2c1d792} /* (0, 26, 24) {real, imag} */,
  {32'h42b4f015, 32'hc107cb40} /* (0, 26, 23) {real, imag} */,
  {32'hc28e4698, 32'hc1522d78} /* (0, 26, 22) {real, imag} */,
  {32'hc2215500, 32'hc23f011b} /* (0, 26, 21) {real, imag} */,
  {32'h41b6bdde, 32'hc11358c8} /* (0, 26, 20) {real, imag} */,
  {32'hbf863dc0, 32'hc1de6f78} /* (0, 26, 19) {real, imag} */,
  {32'hc0073030, 32'hc17d313e} /* (0, 26, 18) {real, imag} */,
  {32'h40a6365c, 32'h40f75e34} /* (0, 26, 17) {real, imag} */,
  {32'hc0868e48, 32'h00000000} /* (0, 26, 16) {real, imag} */,
  {32'h40a6365c, 32'hc0f75e34} /* (0, 26, 15) {real, imag} */,
  {32'hc0073030, 32'h417d313e} /* (0, 26, 14) {real, imag} */,
  {32'hbf863dc0, 32'h41de6f78} /* (0, 26, 13) {real, imag} */,
  {32'h41b6bdde, 32'h411358c8} /* (0, 26, 12) {real, imag} */,
  {32'hc2215500, 32'h423f011b} /* (0, 26, 11) {real, imag} */,
  {32'hc28e4698, 32'h41522d78} /* (0, 26, 10) {real, imag} */,
  {32'h42b4f015, 32'h4107cb40} /* (0, 26, 9) {real, imag} */,
  {32'h4255470a, 32'h42c1d792} /* (0, 26, 8) {real, imag} */,
  {32'h41e0f145, 32'hc28be12f} /* (0, 26, 7) {real, imag} */,
  {32'h41ca84b3, 32'h40a2f3c0} /* (0, 26, 6) {real, imag} */,
  {32'h4311c5c2, 32'h420018cf} /* (0, 26, 5) {real, imag} */,
  {32'hc2fa53e6, 32'hc2e19571} /* (0, 26, 4) {real, imag} */,
  {32'hc212b92c, 32'h4229c27f} /* (0, 26, 3) {real, imag} */,
  {32'h433c427b, 32'hc2aec14d} /* (0, 26, 2) {real, imag} */,
  {32'hc4496816, 32'hc27bd300} /* (0, 26, 1) {real, imag} */,
  {32'hc392af36, 32'h00000000} /* (0, 26, 0) {real, imag} */,
  {32'hc465e3ba, 32'hc3494f78} /* (0, 25, 31) {real, imag} */,
  {32'h438060fb, 32'h4342b451} /* (0, 25, 30) {real, imag} */,
  {32'hc2c0a8f9, 32'h418ad2c8} /* (0, 25, 29) {real, imag} */,
  {32'hc30cdbf4, 32'h41f93a00} /* (0, 25, 28) {real, imag} */,
  {32'h434f5b8a, 32'hc3044082} /* (0, 25, 27) {real, imag} */,
  {32'h42e882e8, 32'hc1881342} /* (0, 25, 26) {real, imag} */,
  {32'hc107bb3e, 32'h42e3efc8} /* (0, 25, 25) {real, imag} */,
  {32'h41c2320d, 32'hc327d723} /* (0, 25, 24) {real, imag} */,
  {32'hc2978c53, 32'hc264e13f} /* (0, 25, 23) {real, imag} */,
  {32'h4219b63f, 32'hc24714e6} /* (0, 25, 22) {real, imag} */,
  {32'hc29254a6, 32'h4195b51c} /* (0, 25, 21) {real, imag} */,
  {32'h41885bec, 32'hc20c42a6} /* (0, 25, 20) {real, imag} */,
  {32'hc143f4c6, 32'hc0fc45b8} /* (0, 25, 19) {real, imag} */,
  {32'hc187c30d, 32'h41203879} /* (0, 25, 18) {real, imag} */,
  {32'hc202d125, 32'hc24d6543} /* (0, 25, 17) {real, imag} */,
  {32'h424ab017, 32'h00000000} /* (0, 25, 16) {real, imag} */,
  {32'hc202d125, 32'h424d6543} /* (0, 25, 15) {real, imag} */,
  {32'hc187c30d, 32'hc1203879} /* (0, 25, 14) {real, imag} */,
  {32'hc143f4c6, 32'h40fc45b8} /* (0, 25, 13) {real, imag} */,
  {32'h41885bec, 32'h420c42a6} /* (0, 25, 12) {real, imag} */,
  {32'hc29254a6, 32'hc195b51c} /* (0, 25, 11) {real, imag} */,
  {32'h4219b63f, 32'h424714e6} /* (0, 25, 10) {real, imag} */,
  {32'hc2978c53, 32'h4264e13f} /* (0, 25, 9) {real, imag} */,
  {32'h41c2320d, 32'h4327d723} /* (0, 25, 8) {real, imag} */,
  {32'hc107bb3e, 32'hc2e3efc8} /* (0, 25, 7) {real, imag} */,
  {32'h42e882e8, 32'h41881342} /* (0, 25, 6) {real, imag} */,
  {32'h434f5b8a, 32'h43044082} /* (0, 25, 5) {real, imag} */,
  {32'hc30cdbf4, 32'hc1f93a00} /* (0, 25, 4) {real, imag} */,
  {32'hc2c0a8f9, 32'hc18ad2c8} /* (0, 25, 3) {real, imag} */,
  {32'h438060fb, 32'hc342b451} /* (0, 25, 2) {real, imag} */,
  {32'hc465e3ba, 32'h43494f78} /* (0, 25, 1) {real, imag} */,
  {32'hc39102c1, 32'h00000000} /* (0, 25, 0) {real, imag} */,
  {32'hc428e684, 32'hc255784c} /* (0, 24, 31) {real, imag} */,
  {32'h433ad7e5, 32'h42b51054} /* (0, 24, 30) {real, imag} */,
  {32'hc1d93086, 32'h41e27866} /* (0, 24, 29) {real, imag} */,
  {32'hc3230d0c, 32'hc206a040} /* (0, 24, 28) {real, imag} */,
  {32'h42cfdd8c, 32'hc2ae7034} /* (0, 24, 27) {real, imag} */,
  {32'hc1d94dbe, 32'h3e191a00} /* (0, 24, 26) {real, imag} */,
  {32'h40b7a2a0, 32'h420fcff4} /* (0, 24, 25) {real, imag} */,
  {32'hc17fe01c, 32'hc19c468e} /* (0, 24, 24) {real, imag} */,
  {32'h4115a7e8, 32'hc28b6822} /* (0, 24, 23) {real, imag} */,
  {32'h4282e808, 32'h42959f62} /* (0, 24, 22) {real, imag} */,
  {32'hc2507fda, 32'hc1676f1e} /* (0, 24, 21) {real, imag} */,
  {32'hc203f76e, 32'h407ef254} /* (0, 24, 20) {real, imag} */,
  {32'hc23d6c31, 32'h417c96da} /* (0, 24, 19) {real, imag} */,
  {32'h42268cf8, 32'hc22e4a31} /* (0, 24, 18) {real, imag} */,
  {32'hc201b96a, 32'h4226f5b3} /* (0, 24, 17) {real, imag} */,
  {32'hc1630497, 32'h00000000} /* (0, 24, 16) {real, imag} */,
  {32'hc201b96a, 32'hc226f5b3} /* (0, 24, 15) {real, imag} */,
  {32'h42268cf8, 32'h422e4a31} /* (0, 24, 14) {real, imag} */,
  {32'hc23d6c31, 32'hc17c96da} /* (0, 24, 13) {real, imag} */,
  {32'hc203f76e, 32'hc07ef254} /* (0, 24, 12) {real, imag} */,
  {32'hc2507fda, 32'h41676f1e} /* (0, 24, 11) {real, imag} */,
  {32'h4282e808, 32'hc2959f62} /* (0, 24, 10) {real, imag} */,
  {32'h4115a7e8, 32'h428b6822} /* (0, 24, 9) {real, imag} */,
  {32'hc17fe01c, 32'h419c468e} /* (0, 24, 8) {real, imag} */,
  {32'h40b7a2a0, 32'hc20fcff4} /* (0, 24, 7) {real, imag} */,
  {32'hc1d94dbe, 32'hbe191a00} /* (0, 24, 6) {real, imag} */,
  {32'h42cfdd8c, 32'h42ae7034} /* (0, 24, 5) {real, imag} */,
  {32'hc3230d0c, 32'h4206a040} /* (0, 24, 4) {real, imag} */,
  {32'hc1d93086, 32'hc1e27866} /* (0, 24, 3) {real, imag} */,
  {32'h433ad7e5, 32'hc2b51054} /* (0, 24, 2) {real, imag} */,
  {32'hc428e684, 32'h4255784c} /* (0, 24, 1) {real, imag} */,
  {32'hc2442210, 32'h00000000} /* (0, 24, 0) {real, imag} */,
  {32'hc4149373, 32'h424a0f22} /* (0, 23, 31) {real, imag} */,
  {32'h42b3c324, 32'h42e6bf66} /* (0, 23, 30) {real, imag} */,
  {32'h42dc5787, 32'h4205e1d4} /* (0, 23, 29) {real, imag} */,
  {32'hc282d814, 32'hc17d6156} /* (0, 23, 28) {real, imag} */,
  {32'h42d8faec, 32'hc27423aa} /* (0, 23, 27) {real, imag} */,
  {32'hc214eae2, 32'hc12a94a1} /* (0, 23, 26) {real, imag} */,
  {32'hc279b577, 32'h4266087d} /* (0, 23, 25) {real, imag} */,
  {32'h428e1f99, 32'h411417a0} /* (0, 23, 24) {real, imag} */,
  {32'hc13b846e, 32'hc1e57dbf} /* (0, 23, 23) {real, imag} */,
  {32'hc1913fd4, 32'hc203a6f1} /* (0, 23, 22) {real, imag} */,
  {32'h4265c1c5, 32'hc1a34e38} /* (0, 23, 21) {real, imag} */,
  {32'h41aa2ea1, 32'h411787fc} /* (0, 23, 20) {real, imag} */,
  {32'h41174272, 32'h40a3bca2} /* (0, 23, 19) {real, imag} */,
  {32'h420872b5, 32'hc2095eb8} /* (0, 23, 18) {real, imag} */,
  {32'hc267c1ea, 32'hc1f6d19b} /* (0, 23, 17) {real, imag} */,
  {32'hc22155db, 32'h00000000} /* (0, 23, 16) {real, imag} */,
  {32'hc267c1ea, 32'h41f6d19b} /* (0, 23, 15) {real, imag} */,
  {32'h420872b5, 32'h42095eb8} /* (0, 23, 14) {real, imag} */,
  {32'h41174272, 32'hc0a3bca2} /* (0, 23, 13) {real, imag} */,
  {32'h41aa2ea1, 32'hc11787fc} /* (0, 23, 12) {real, imag} */,
  {32'h4265c1c5, 32'h41a34e38} /* (0, 23, 11) {real, imag} */,
  {32'hc1913fd4, 32'h4203a6f1} /* (0, 23, 10) {real, imag} */,
  {32'hc13b846e, 32'h41e57dbf} /* (0, 23, 9) {real, imag} */,
  {32'h428e1f99, 32'hc11417a0} /* (0, 23, 8) {real, imag} */,
  {32'hc279b577, 32'hc266087d} /* (0, 23, 7) {real, imag} */,
  {32'hc214eae2, 32'h412a94a1} /* (0, 23, 6) {real, imag} */,
  {32'h42d8faec, 32'h427423aa} /* (0, 23, 5) {real, imag} */,
  {32'hc282d814, 32'h417d6156} /* (0, 23, 4) {real, imag} */,
  {32'h42dc5787, 32'hc205e1d4} /* (0, 23, 3) {real, imag} */,
  {32'h42b3c324, 32'hc2e6bf66} /* (0, 23, 2) {real, imag} */,
  {32'hc4149373, 32'hc24a0f22} /* (0, 23, 1) {real, imag} */,
  {32'hc041d100, 32'h00000000} /* (0, 23, 0) {real, imag} */,
  {32'hc3f7a3d4, 32'h43139836} /* (0, 22, 31) {real, imag} */,
  {32'h42e44362, 32'h4220c64e} /* (0, 22, 30) {real, imag} */,
  {32'h43170bca, 32'h429c06ca} /* (0, 22, 29) {real, imag} */,
  {32'hc2d55b81, 32'hc23660b9} /* (0, 22, 28) {real, imag} */,
  {32'h42c9833b, 32'hc2a29d9a} /* (0, 22, 27) {real, imag} */,
  {32'hc1eec9ac, 32'hc08c1b1c} /* (0, 22, 26) {real, imag} */,
  {32'hc2d00e68, 32'hc0ecb3a0} /* (0, 22, 25) {real, imag} */,
  {32'h426d69b8, 32'hc027cc86} /* (0, 22, 24) {real, imag} */,
  {32'hc19ead3d, 32'h416b227a} /* (0, 22, 23) {real, imag} */,
  {32'h42274051, 32'hc10aa346} /* (0, 22, 22) {real, imag} */,
  {32'hc193aba9, 32'h417f7860} /* (0, 22, 21) {real, imag} */,
  {32'h4248c54b, 32'hc18e64d1} /* (0, 22, 20) {real, imag} */,
  {32'hc0071f54, 32'h429b18de} /* (0, 22, 19) {real, imag} */,
  {32'hc2526b2a, 32'h41fc5ad2} /* (0, 22, 18) {real, imag} */,
  {32'h3e593bc0, 32'h41b3f14c} /* (0, 22, 17) {real, imag} */,
  {32'hc24cbe82, 32'h00000000} /* (0, 22, 16) {real, imag} */,
  {32'h3e593bc0, 32'hc1b3f14c} /* (0, 22, 15) {real, imag} */,
  {32'hc2526b2a, 32'hc1fc5ad2} /* (0, 22, 14) {real, imag} */,
  {32'hc0071f54, 32'hc29b18de} /* (0, 22, 13) {real, imag} */,
  {32'h4248c54b, 32'h418e64d1} /* (0, 22, 12) {real, imag} */,
  {32'hc193aba9, 32'hc17f7860} /* (0, 22, 11) {real, imag} */,
  {32'h42274051, 32'h410aa346} /* (0, 22, 10) {real, imag} */,
  {32'hc19ead3d, 32'hc16b227a} /* (0, 22, 9) {real, imag} */,
  {32'h426d69b8, 32'h4027cc86} /* (0, 22, 8) {real, imag} */,
  {32'hc2d00e68, 32'h40ecb3a0} /* (0, 22, 7) {real, imag} */,
  {32'hc1eec9ac, 32'h408c1b1c} /* (0, 22, 6) {real, imag} */,
  {32'h42c9833b, 32'h42a29d9a} /* (0, 22, 5) {real, imag} */,
  {32'hc2d55b81, 32'h423660b9} /* (0, 22, 4) {real, imag} */,
  {32'h43170bca, 32'hc29c06ca} /* (0, 22, 3) {real, imag} */,
  {32'h42e44362, 32'hc220c64e} /* (0, 22, 2) {real, imag} */,
  {32'hc3f7a3d4, 32'hc3139836} /* (0, 22, 1) {real, imag} */,
  {32'hc0968080, 32'h00000000} /* (0, 22, 0) {real, imag} */,
  {32'hc38a8924, 32'h42cc8096} /* (0, 21, 31) {real, imag} */,
  {32'h40303e40, 32'h41ad55b6} /* (0, 21, 30) {real, imag} */,
  {32'h4285aa18, 32'h42cbd848} /* (0, 21, 29) {real, imag} */,
  {32'hc2701e51, 32'hc178b690} /* (0, 21, 28) {real, imag} */,
  {32'h4206af79, 32'hc2854b02} /* (0, 21, 27) {real, imag} */,
  {32'hc24a0881, 32'h418a9ebf} /* (0, 21, 26) {real, imag} */,
  {32'hc1be8666, 32'hc302c042} /* (0, 21, 25) {real, imag} */,
  {32'hc21e7927, 32'h4142dc50} /* (0, 21, 24) {real, imag} */,
  {32'hc18e4e97, 32'h42b636f6} /* (0, 21, 23) {real, imag} */,
  {32'hc0092208, 32'h4237d58f} /* (0, 21, 22) {real, imag} */,
  {32'h4212ced0, 32'hc269cc9a} /* (0, 21, 21) {real, imag} */,
  {32'h4288acbf, 32'hc2304856} /* (0, 21, 20) {real, imag} */,
  {32'hc08af83a, 32'h41eefe02} /* (0, 21, 19) {real, imag} */,
  {32'hc1de1ba8, 32'hc2a01f1c} /* (0, 21, 18) {real, imag} */,
  {32'h41008ca6, 32'hc19abcb8} /* (0, 21, 17) {real, imag} */,
  {32'hc1a0d4df, 32'h00000000} /* (0, 21, 16) {real, imag} */,
  {32'h41008ca6, 32'h419abcb8} /* (0, 21, 15) {real, imag} */,
  {32'hc1de1ba8, 32'h42a01f1c} /* (0, 21, 14) {real, imag} */,
  {32'hc08af83a, 32'hc1eefe02} /* (0, 21, 13) {real, imag} */,
  {32'h4288acbf, 32'h42304856} /* (0, 21, 12) {real, imag} */,
  {32'h4212ced0, 32'h4269cc9a} /* (0, 21, 11) {real, imag} */,
  {32'hc0092208, 32'hc237d58f} /* (0, 21, 10) {real, imag} */,
  {32'hc18e4e97, 32'hc2b636f6} /* (0, 21, 9) {real, imag} */,
  {32'hc21e7927, 32'hc142dc50} /* (0, 21, 8) {real, imag} */,
  {32'hc1be8666, 32'h4302c042} /* (0, 21, 7) {real, imag} */,
  {32'hc24a0881, 32'hc18a9ebf} /* (0, 21, 6) {real, imag} */,
  {32'h4206af79, 32'h42854b02} /* (0, 21, 5) {real, imag} */,
  {32'hc2701e51, 32'h4178b690} /* (0, 21, 4) {real, imag} */,
  {32'h4285aa18, 32'hc2cbd848} /* (0, 21, 3) {real, imag} */,
  {32'h40303e40, 32'hc1ad55b6} /* (0, 21, 2) {real, imag} */,
  {32'hc38a8924, 32'hc2cc8096} /* (0, 21, 1) {real, imag} */,
  {32'h41c72f00, 32'h00000000} /* (0, 21, 0) {real, imag} */,
  {32'h42d86d78, 32'hc2aea494} /* (0, 20, 31) {real, imag} */,
  {32'hc376523f, 32'h41b3d514} /* (0, 20, 30) {real, imag} */,
  {32'hc2336daf, 32'h42e9b033} /* (0, 20, 29) {real, imag} */,
  {32'h42273987, 32'hc201f5cb} /* (0, 20, 28) {real, imag} */,
  {32'hc20a2e2e, 32'hc2b98f28} /* (0, 20, 27) {real, imag} */,
  {32'hc1c6ff2e, 32'h425d654a} /* (0, 20, 26) {real, imag} */,
  {32'hc2a34d31, 32'hc237cd54} /* (0, 20, 25) {real, imag} */,
  {32'h421b988b, 32'h42213af0} /* (0, 20, 24) {real, imag} */,
  {32'h41ecdee5, 32'h40547320} /* (0, 20, 23) {real, imag} */,
  {32'hc2091f60, 32'hc24f401f} /* (0, 20, 22) {real, imag} */,
  {32'h419a618b, 32'h41da8d1a} /* (0, 20, 21) {real, imag} */,
  {32'h42637d6d, 32'h419b04c4} /* (0, 20, 20) {real, imag} */,
  {32'hc285ffa4, 32'hc1235a88} /* (0, 20, 19) {real, imag} */,
  {32'h4257fdb0, 32'hc22a86a0} /* (0, 20, 18) {real, imag} */,
  {32'hc20e46d1, 32'hc1d5241c} /* (0, 20, 17) {real, imag} */,
  {32'h41a19b74, 32'h00000000} /* (0, 20, 16) {real, imag} */,
  {32'hc20e46d1, 32'h41d5241c} /* (0, 20, 15) {real, imag} */,
  {32'h4257fdb0, 32'h422a86a0} /* (0, 20, 14) {real, imag} */,
  {32'hc285ffa4, 32'h41235a88} /* (0, 20, 13) {real, imag} */,
  {32'h42637d6d, 32'hc19b04c4} /* (0, 20, 12) {real, imag} */,
  {32'h419a618b, 32'hc1da8d1a} /* (0, 20, 11) {real, imag} */,
  {32'hc2091f60, 32'h424f401f} /* (0, 20, 10) {real, imag} */,
  {32'h41ecdee5, 32'hc0547320} /* (0, 20, 9) {real, imag} */,
  {32'h421b988b, 32'hc2213af0} /* (0, 20, 8) {real, imag} */,
  {32'hc2a34d31, 32'h4237cd54} /* (0, 20, 7) {real, imag} */,
  {32'hc1c6ff2e, 32'hc25d654a} /* (0, 20, 6) {real, imag} */,
  {32'hc20a2e2e, 32'h42b98f28} /* (0, 20, 5) {real, imag} */,
  {32'h42273987, 32'h4201f5cb} /* (0, 20, 4) {real, imag} */,
  {32'hc2336daf, 32'hc2e9b033} /* (0, 20, 3) {real, imag} */,
  {32'hc376523f, 32'hc1b3d514} /* (0, 20, 2) {real, imag} */,
  {32'h42d86d78, 32'h42aea494} /* (0, 20, 1) {real, imag} */,
  {32'h4399354e, 32'h00000000} /* (0, 20, 0) {real, imag} */,
  {32'h43930610, 32'hc2e121fc} /* (0, 19, 31) {real, imag} */,
  {32'hc35c738b, 32'h413891c8} /* (0, 19, 30) {real, imag} */,
  {32'hc273aed3, 32'h42033c96} /* (0, 19, 29) {real, imag} */,
  {32'hc0f3e798, 32'hc28d94d6} /* (0, 19, 28) {real, imag} */,
  {32'h3f80e400, 32'hc0bed990} /* (0, 19, 27) {real, imag} */,
  {32'hc290d589, 32'hc28bddf2} /* (0, 19, 26) {real, imag} */,
  {32'hc216eb00, 32'hc23ada10} /* (0, 19, 25) {real, imag} */,
  {32'h41425f56, 32'h42a1f3d4} /* (0, 19, 24) {real, imag} */,
  {32'hc20346cc, 32'h4191d3ca} /* (0, 19, 23) {real, imag} */,
  {32'h419d9e80, 32'h42275e2b} /* (0, 19, 22) {real, imag} */,
  {32'hc20491c6, 32'h42e27822} /* (0, 19, 21) {real, imag} */,
  {32'hc22116e8, 32'h4135e7d8} /* (0, 19, 20) {real, imag} */,
  {32'h41af05f7, 32'hc1201752} /* (0, 19, 19) {real, imag} */,
  {32'h41df83b4, 32'hc01b0902} /* (0, 19, 18) {real, imag} */,
  {32'h41202915, 32'h4002dbec} /* (0, 19, 17) {real, imag} */,
  {32'hc13943fc, 32'h00000000} /* (0, 19, 16) {real, imag} */,
  {32'h41202915, 32'hc002dbec} /* (0, 19, 15) {real, imag} */,
  {32'h41df83b4, 32'h401b0902} /* (0, 19, 14) {real, imag} */,
  {32'h41af05f7, 32'h41201752} /* (0, 19, 13) {real, imag} */,
  {32'hc22116e8, 32'hc135e7d8} /* (0, 19, 12) {real, imag} */,
  {32'hc20491c6, 32'hc2e27822} /* (0, 19, 11) {real, imag} */,
  {32'h419d9e80, 32'hc2275e2b} /* (0, 19, 10) {real, imag} */,
  {32'hc20346cc, 32'hc191d3ca} /* (0, 19, 9) {real, imag} */,
  {32'h41425f56, 32'hc2a1f3d4} /* (0, 19, 8) {real, imag} */,
  {32'hc216eb00, 32'h423ada10} /* (0, 19, 7) {real, imag} */,
  {32'hc290d589, 32'h428bddf2} /* (0, 19, 6) {real, imag} */,
  {32'h3f80e400, 32'h40bed990} /* (0, 19, 5) {real, imag} */,
  {32'hc0f3e798, 32'h428d94d6} /* (0, 19, 4) {real, imag} */,
  {32'hc273aed3, 32'hc2033c96} /* (0, 19, 3) {real, imag} */,
  {32'hc35c738b, 32'hc13891c8} /* (0, 19, 2) {real, imag} */,
  {32'h43930610, 32'h42e121fc} /* (0, 19, 1) {real, imag} */,
  {32'h43fa9a1e, 32'h00000000} /* (0, 19, 0) {real, imag} */,
  {32'h43d59edf, 32'hc327a5de} /* (0, 18, 31) {real, imag} */,
  {32'hc3916d98, 32'h42fc2471} /* (0, 18, 30) {real, imag} */,
  {32'hc2cd0ad0, 32'h42724364} /* (0, 18, 29) {real, imag} */,
  {32'h42c0e467, 32'hc2b3d5cb} /* (0, 18, 28) {real, imag} */,
  {32'hc27b866e, 32'h41865d4d} /* (0, 18, 27) {real, imag} */,
  {32'hc0e7f62e, 32'hc28add85} /* (0, 18, 26) {real, imag} */,
  {32'hc27a7e24, 32'h42bfd66a} /* (0, 18, 25) {real, imag} */,
  {32'hc20e2ba7, 32'hc1a66d03} /* (0, 18, 24) {real, imag} */,
  {32'hc204f41d, 32'h4116e61c} /* (0, 18, 23) {real, imag} */,
  {32'hc1f1107c, 32'h424e7f31} /* (0, 18, 22) {real, imag} */,
  {32'hc10d4245, 32'h41f76682} /* (0, 18, 21) {real, imag} */,
  {32'h41fac042, 32'hc20bc3e8} /* (0, 18, 20) {real, imag} */,
  {32'hc22137a8, 32'hc1833210} /* (0, 18, 19) {real, imag} */,
  {32'hc21dc45f, 32'h423784a4} /* (0, 18, 18) {real, imag} */,
  {32'hc215800c, 32'h412834b0} /* (0, 18, 17) {real, imag} */,
  {32'h3f9f5f95, 32'h00000000} /* (0, 18, 16) {real, imag} */,
  {32'hc215800c, 32'hc12834b0} /* (0, 18, 15) {real, imag} */,
  {32'hc21dc45f, 32'hc23784a4} /* (0, 18, 14) {real, imag} */,
  {32'hc22137a8, 32'h41833210} /* (0, 18, 13) {real, imag} */,
  {32'h41fac042, 32'h420bc3e8} /* (0, 18, 12) {real, imag} */,
  {32'hc10d4245, 32'hc1f76682} /* (0, 18, 11) {real, imag} */,
  {32'hc1f1107c, 32'hc24e7f31} /* (0, 18, 10) {real, imag} */,
  {32'hc204f41d, 32'hc116e61c} /* (0, 18, 9) {real, imag} */,
  {32'hc20e2ba7, 32'h41a66d03} /* (0, 18, 8) {real, imag} */,
  {32'hc27a7e24, 32'hc2bfd66a} /* (0, 18, 7) {real, imag} */,
  {32'hc0e7f62e, 32'h428add85} /* (0, 18, 6) {real, imag} */,
  {32'hc27b866e, 32'hc1865d4d} /* (0, 18, 5) {real, imag} */,
  {32'h42c0e467, 32'h42b3d5cb} /* (0, 18, 4) {real, imag} */,
  {32'hc2cd0ad0, 32'hc2724364} /* (0, 18, 3) {real, imag} */,
  {32'hc3916d98, 32'hc2fc2471} /* (0, 18, 2) {real, imag} */,
  {32'h43d59edf, 32'h4327a5de} /* (0, 18, 1) {real, imag} */,
  {32'h43d00180, 32'h00000000} /* (0, 18, 0) {real, imag} */,
  {32'h43cfe619, 32'hc344ede8} /* (0, 17, 31) {real, imag} */,
  {32'hc3b45ad0, 32'hc182ee14} /* (0, 17, 30) {real, imag} */,
  {32'hc1725cdc, 32'hc1997124} /* (0, 17, 29) {real, imag} */,
  {32'h42358aaf, 32'hc1b1c08e} /* (0, 17, 28) {real, imag} */,
  {32'hbf10cc00, 32'h4278c733} /* (0, 17, 27) {real, imag} */,
  {32'h41aa6e61, 32'hc2292b4c} /* (0, 17, 26) {real, imag} */,
  {32'h4190e5be, 32'h427fe156} /* (0, 17, 25) {real, imag} */,
  {32'hc1095478, 32'h400c1370} /* (0, 17, 24) {real, imag} */,
  {32'h40f45068, 32'hc20d999e} /* (0, 17, 23) {real, imag} */,
  {32'h428d8486, 32'hc1417cee} /* (0, 17, 22) {real, imag} */,
  {32'hc2b1e4d3, 32'h41fbf8a8} /* (0, 17, 21) {real, imag} */,
  {32'h41abf3bb, 32'h40e49f70} /* (0, 17, 20) {real, imag} */,
  {32'hc212e14a, 32'hc123a052} /* (0, 17, 19) {real, imag} */,
  {32'hc09c5890, 32'h42318469} /* (0, 17, 18) {real, imag} */,
  {32'hc0592322, 32'h4156db13} /* (0, 17, 17) {real, imag} */,
  {32'h42215d93, 32'h00000000} /* (0, 17, 16) {real, imag} */,
  {32'hc0592322, 32'hc156db13} /* (0, 17, 15) {real, imag} */,
  {32'hc09c5890, 32'hc2318469} /* (0, 17, 14) {real, imag} */,
  {32'hc212e14a, 32'h4123a052} /* (0, 17, 13) {real, imag} */,
  {32'h41abf3bb, 32'hc0e49f70} /* (0, 17, 12) {real, imag} */,
  {32'hc2b1e4d3, 32'hc1fbf8a8} /* (0, 17, 11) {real, imag} */,
  {32'h428d8486, 32'h41417cee} /* (0, 17, 10) {real, imag} */,
  {32'h40f45068, 32'h420d999e} /* (0, 17, 9) {real, imag} */,
  {32'hc1095478, 32'hc00c1370} /* (0, 17, 8) {real, imag} */,
  {32'h4190e5be, 32'hc27fe156} /* (0, 17, 7) {real, imag} */,
  {32'h41aa6e61, 32'h42292b4c} /* (0, 17, 6) {real, imag} */,
  {32'hbf10cc00, 32'hc278c733} /* (0, 17, 5) {real, imag} */,
  {32'h42358aaf, 32'h41b1c08e} /* (0, 17, 4) {real, imag} */,
  {32'hc1725cdc, 32'h41997124} /* (0, 17, 3) {real, imag} */,
  {32'hc3b45ad0, 32'h4182ee14} /* (0, 17, 2) {real, imag} */,
  {32'h43cfe619, 32'h4344ede8} /* (0, 17, 1) {real, imag} */,
  {32'h43d0829d, 32'h00000000} /* (0, 17, 0) {real, imag} */,
  {32'h43ff9562, 32'hc3353312} /* (0, 16, 31) {real, imag} */,
  {32'hc3e303b1, 32'h414d824e} /* (0, 16, 30) {real, imag} */,
  {32'hc207b097, 32'hc35a41a8} /* (0, 16, 29) {real, imag} */,
  {32'h42b6ae6a, 32'h41446fb8} /* (0, 16, 28) {real, imag} */,
  {32'hc28da400, 32'h43046e1b} /* (0, 16, 27) {real, imag} */,
  {32'hc211b5a4, 32'hc18a8da8} /* (0, 16, 26) {real, imag} */,
  {32'h429de84d, 32'h41cbab40} /* (0, 16, 25) {real, imag} */,
  {32'hc2526bac, 32'h422be942} /* (0, 16, 24) {real, imag} */,
  {32'h41a2604d, 32'h42171b0b} /* (0, 16, 23) {real, imag} */,
  {32'hc00ed288, 32'hc2711194} /* (0, 16, 22) {real, imag} */,
  {32'h41edf9d5, 32'h422af2ec} /* (0, 16, 21) {real, imag} */,
  {32'h415dd7e9, 32'h42a031b5} /* (0, 16, 20) {real, imag} */,
  {32'h410447f4, 32'h41270580} /* (0, 16, 19) {real, imag} */,
  {32'h4273030a, 32'hc2740036} /* (0, 16, 18) {real, imag} */,
  {32'hc1b004dc, 32'h420d669b} /* (0, 16, 17) {real, imag} */,
  {32'h418564a1, 32'h00000000} /* (0, 16, 16) {real, imag} */,
  {32'hc1b004dc, 32'hc20d669b} /* (0, 16, 15) {real, imag} */,
  {32'h4273030a, 32'h42740036} /* (0, 16, 14) {real, imag} */,
  {32'h410447f4, 32'hc1270580} /* (0, 16, 13) {real, imag} */,
  {32'h415dd7e9, 32'hc2a031b5} /* (0, 16, 12) {real, imag} */,
  {32'h41edf9d5, 32'hc22af2ec} /* (0, 16, 11) {real, imag} */,
  {32'hc00ed288, 32'h42711194} /* (0, 16, 10) {real, imag} */,
  {32'h41a2604d, 32'hc2171b0b} /* (0, 16, 9) {real, imag} */,
  {32'hc2526bac, 32'hc22be942} /* (0, 16, 8) {real, imag} */,
  {32'h429de84d, 32'hc1cbab40} /* (0, 16, 7) {real, imag} */,
  {32'hc211b5a4, 32'h418a8da8} /* (0, 16, 6) {real, imag} */,
  {32'hc28da400, 32'hc3046e1b} /* (0, 16, 5) {real, imag} */,
  {32'h42b6ae6a, 32'hc1446fb8} /* (0, 16, 4) {real, imag} */,
  {32'hc207b097, 32'h435a41a8} /* (0, 16, 3) {real, imag} */,
  {32'hc3e303b1, 32'hc14d824e} /* (0, 16, 2) {real, imag} */,
  {32'h43ff9562, 32'h43353312} /* (0, 16, 1) {real, imag} */,
  {32'h440487c7, 32'h00000000} /* (0, 16, 0) {real, imag} */,
  {32'h44346e38, 32'hc36629d8} /* (0, 15, 31) {real, imag} */,
  {32'hc36241c8, 32'h43690fde} /* (0, 15, 30) {real, imag} */,
  {32'hc2fd9cbc, 32'hc300145c} /* (0, 15, 29) {real, imag} */,
  {32'h422bcd99, 32'h41285800} /* (0, 15, 28) {real, imag} */,
  {32'hc2fadce1, 32'h4289b428} /* (0, 15, 27) {real, imag} */,
  {32'h41b04047, 32'hc1d46bb8} /* (0, 15, 26) {real, imag} */,
  {32'h4211d716, 32'h4283a84f} /* (0, 15, 25) {real, imag} */,
  {32'hc2a32795, 32'h427e69c5} /* (0, 15, 24) {real, imag} */,
  {32'hc27a939d, 32'hc2552158} /* (0, 15, 23) {real, imag} */,
  {32'h4135b25c, 32'h42096540} /* (0, 15, 22) {real, imag} */,
  {32'hc196f2b4, 32'hc1ad0bd4} /* (0, 15, 21) {real, imag} */,
  {32'hc1dc7e5d, 32'hc142983c} /* (0, 15, 20) {real, imag} */,
  {32'hc2a6e389, 32'hc1ffcccf} /* (0, 15, 19) {real, imag} */,
  {32'h4185c13d, 32'hc290b172} /* (0, 15, 18) {real, imag} */,
  {32'h4096a1a1, 32'hc1a61e3a} /* (0, 15, 17) {real, imag} */,
  {32'hc1e3b9f2, 32'h00000000} /* (0, 15, 16) {real, imag} */,
  {32'h4096a1a1, 32'h41a61e3a} /* (0, 15, 15) {real, imag} */,
  {32'h4185c13d, 32'h4290b172} /* (0, 15, 14) {real, imag} */,
  {32'hc2a6e389, 32'h41ffcccf} /* (0, 15, 13) {real, imag} */,
  {32'hc1dc7e5d, 32'h4142983c} /* (0, 15, 12) {real, imag} */,
  {32'hc196f2b4, 32'h41ad0bd4} /* (0, 15, 11) {real, imag} */,
  {32'h4135b25c, 32'hc2096540} /* (0, 15, 10) {real, imag} */,
  {32'hc27a939d, 32'h42552158} /* (0, 15, 9) {real, imag} */,
  {32'hc2a32795, 32'hc27e69c5} /* (0, 15, 8) {real, imag} */,
  {32'h4211d716, 32'hc283a84f} /* (0, 15, 7) {real, imag} */,
  {32'h41b04047, 32'h41d46bb8} /* (0, 15, 6) {real, imag} */,
  {32'hc2fadce1, 32'hc289b428} /* (0, 15, 5) {real, imag} */,
  {32'h422bcd99, 32'hc1285800} /* (0, 15, 4) {real, imag} */,
  {32'hc2fd9cbc, 32'h4300145c} /* (0, 15, 3) {real, imag} */,
  {32'hc36241c8, 32'hc3690fde} /* (0, 15, 2) {real, imag} */,
  {32'h44346e38, 32'h436629d8} /* (0, 15, 1) {real, imag} */,
  {32'h43941f2b, 32'h00000000} /* (0, 15, 0) {real, imag} */,
  {32'h442bd902, 32'hc318296e} /* (0, 14, 31) {real, imag} */,
  {32'hc354b40e, 32'h42a4c60f} /* (0, 14, 30) {real, imag} */,
  {32'hc2a9169e, 32'h42b876c4} /* (0, 14, 29) {real, imag} */,
  {32'hc1fc8244, 32'hc211aa18} /* (0, 14, 28) {real, imag} */,
  {32'hc2a0a341, 32'h428e2c1b} /* (0, 14, 27) {real, imag} */,
  {32'h40fe4642, 32'hc2007fe6} /* (0, 14, 26) {real, imag} */,
  {32'h4210b898, 32'h4111dfe8} /* (0, 14, 25) {real, imag} */,
  {32'hc13c2cbc, 32'hc0d49944} /* (0, 14, 24) {real, imag} */,
  {32'hbea36680, 32'h4251504a} /* (0, 14, 23) {real, imag} */,
  {32'h4190e45a, 32'hbf802da0} /* (0, 14, 22) {real, imag} */,
  {32'hc20a4927, 32'hc12a59cc} /* (0, 14, 21) {real, imag} */,
  {32'h42139931, 32'hc224ff16} /* (0, 14, 20) {real, imag} */,
  {32'hc1eb5ba0, 32'h41bf2b02} /* (0, 14, 19) {real, imag} */,
  {32'h4209f7e1, 32'h41ca6b28} /* (0, 14, 18) {real, imag} */,
  {32'hc14336c6, 32'h40848e9c} /* (0, 14, 17) {real, imag} */,
  {32'hbe2bb358, 32'h00000000} /* (0, 14, 16) {real, imag} */,
  {32'hc14336c6, 32'hc0848e9c} /* (0, 14, 15) {real, imag} */,
  {32'h4209f7e1, 32'hc1ca6b28} /* (0, 14, 14) {real, imag} */,
  {32'hc1eb5ba0, 32'hc1bf2b02} /* (0, 14, 13) {real, imag} */,
  {32'h42139931, 32'h4224ff16} /* (0, 14, 12) {real, imag} */,
  {32'hc20a4927, 32'h412a59cc} /* (0, 14, 11) {real, imag} */,
  {32'h4190e45a, 32'h3f802da0} /* (0, 14, 10) {real, imag} */,
  {32'hbea36680, 32'hc251504a} /* (0, 14, 9) {real, imag} */,
  {32'hc13c2cbc, 32'h40d49944} /* (0, 14, 8) {real, imag} */,
  {32'h4210b898, 32'hc111dfe8} /* (0, 14, 7) {real, imag} */,
  {32'h40fe4642, 32'h42007fe6} /* (0, 14, 6) {real, imag} */,
  {32'hc2a0a341, 32'hc28e2c1b} /* (0, 14, 5) {real, imag} */,
  {32'hc1fc8244, 32'h4211aa18} /* (0, 14, 4) {real, imag} */,
  {32'hc2a9169e, 32'hc2b876c4} /* (0, 14, 3) {real, imag} */,
  {32'hc354b40e, 32'hc2a4c60f} /* (0, 14, 2) {real, imag} */,
  {32'h442bd902, 32'h4318296e} /* (0, 14, 1) {real, imag} */,
  {32'h43819e2c, 32'h00000000} /* (0, 14, 0) {real, imag} */,
  {32'h442afca0, 32'hc3045110} /* (0, 13, 31) {real, imag} */,
  {32'hc375592d, 32'hc10e08c8} /* (0, 13, 30) {real, imag} */,
  {32'hc2bac1a0, 32'h42aef856} /* (0, 13, 29) {real, imag} */,
  {32'h42953186, 32'hc2c61ea6} /* (0, 13, 28) {real, imag} */,
  {32'hc1f884bc, 32'h42e556e3} /* (0, 13, 27) {real, imag} */,
  {32'hc1e2c599, 32'h426805fc} /* (0, 13, 26) {real, imag} */,
  {32'hc157b8fc, 32'hc136f330} /* (0, 13, 25) {real, imag} */,
  {32'hc26b9362, 32'h4023c250} /* (0, 13, 24) {real, imag} */,
  {32'h42238e22, 32'h4289bc62} /* (0, 13, 23) {real, imag} */,
  {32'h41fe5340, 32'h41142254} /* (0, 13, 22) {real, imag} */,
  {32'hc22fd8ba, 32'h4100e84c} /* (0, 13, 21) {real, imag} */,
  {32'hc12cbf45, 32'h423f5c16} /* (0, 13, 20) {real, imag} */,
  {32'h419836cd, 32'hc22fead0} /* (0, 13, 19) {real, imag} */,
  {32'h4102b405, 32'hc0b64d29} /* (0, 13, 18) {real, imag} */,
  {32'hc12a7797, 32'h41eebac4} /* (0, 13, 17) {real, imag} */,
  {32'hc2569639, 32'h00000000} /* (0, 13, 16) {real, imag} */,
  {32'hc12a7797, 32'hc1eebac4} /* (0, 13, 15) {real, imag} */,
  {32'h4102b405, 32'h40b64d29} /* (0, 13, 14) {real, imag} */,
  {32'h419836cd, 32'h422fead0} /* (0, 13, 13) {real, imag} */,
  {32'hc12cbf45, 32'hc23f5c16} /* (0, 13, 12) {real, imag} */,
  {32'hc22fd8ba, 32'hc100e84c} /* (0, 13, 11) {real, imag} */,
  {32'h41fe5340, 32'hc1142254} /* (0, 13, 10) {real, imag} */,
  {32'h42238e22, 32'hc289bc62} /* (0, 13, 9) {real, imag} */,
  {32'hc26b9362, 32'hc023c250} /* (0, 13, 8) {real, imag} */,
  {32'hc157b8fc, 32'h4136f330} /* (0, 13, 7) {real, imag} */,
  {32'hc1e2c599, 32'hc26805fc} /* (0, 13, 6) {real, imag} */,
  {32'hc1f884bc, 32'hc2e556e3} /* (0, 13, 5) {real, imag} */,
  {32'h42953186, 32'h42c61ea6} /* (0, 13, 4) {real, imag} */,
  {32'hc2bac1a0, 32'hc2aef856} /* (0, 13, 3) {real, imag} */,
  {32'hc375592d, 32'h410e08c8} /* (0, 13, 2) {real, imag} */,
  {32'h442afca0, 32'h43045110} /* (0, 13, 1) {real, imag} */,
  {32'h43477f6b, 32'h00000000} /* (0, 13, 0) {real, imag} */,
  {32'h4405d1ff, 32'hc2fee4dc} /* (0, 12, 31) {real, imag} */,
  {32'hc35eed75, 32'h428da948} /* (0, 12, 30) {real, imag} */,
  {32'hc228a15b, 32'h419d63c4} /* (0, 12, 29) {real, imag} */,
  {32'h41aaf036, 32'hc2cba6e2} /* (0, 12, 28) {real, imag} */,
  {32'h41ee1560, 32'h426d6d1c} /* (0, 12, 27) {real, imag} */,
  {32'h4210435b, 32'h42084c9a} /* (0, 12, 26) {real, imag} */,
  {32'hc15ff468, 32'h400725b8} /* (0, 12, 25) {real, imag} */,
  {32'hc1acf29e, 32'h41ee23a1} /* (0, 12, 24) {real, imag} */,
  {32'h42260008, 32'h41c16a00} /* (0, 12, 23) {real, imag} */,
  {32'hc2b18909, 32'h4121b77c} /* (0, 12, 22) {real, imag} */,
  {32'hc212fbca, 32'h421389d5} /* (0, 12, 21) {real, imag} */,
  {32'hc2b2a0d0, 32'hc12c9183} /* (0, 12, 20) {real, imag} */,
  {32'h41a4c6de, 32'h41bee5ec} /* (0, 12, 19) {real, imag} */,
  {32'hc2018664, 32'h420a18fc} /* (0, 12, 18) {real, imag} */,
  {32'h422ccfcf, 32'h411bddac} /* (0, 12, 17) {real, imag} */,
  {32'hc1ecb6c2, 32'h00000000} /* (0, 12, 16) {real, imag} */,
  {32'h422ccfcf, 32'hc11bddac} /* (0, 12, 15) {real, imag} */,
  {32'hc2018664, 32'hc20a18fc} /* (0, 12, 14) {real, imag} */,
  {32'h41a4c6de, 32'hc1bee5ec} /* (0, 12, 13) {real, imag} */,
  {32'hc2b2a0d0, 32'h412c9183} /* (0, 12, 12) {real, imag} */,
  {32'hc212fbca, 32'hc21389d5} /* (0, 12, 11) {real, imag} */,
  {32'hc2b18909, 32'hc121b77c} /* (0, 12, 10) {real, imag} */,
  {32'h42260008, 32'hc1c16a00} /* (0, 12, 9) {real, imag} */,
  {32'hc1acf29e, 32'hc1ee23a1} /* (0, 12, 8) {real, imag} */,
  {32'hc15ff468, 32'hc00725b8} /* (0, 12, 7) {real, imag} */,
  {32'h4210435b, 32'hc2084c9a} /* (0, 12, 6) {real, imag} */,
  {32'h41ee1560, 32'hc26d6d1c} /* (0, 12, 5) {real, imag} */,
  {32'h41aaf036, 32'h42cba6e2} /* (0, 12, 4) {real, imag} */,
  {32'hc228a15b, 32'hc19d63c4} /* (0, 12, 3) {real, imag} */,
  {32'hc35eed75, 32'hc28da948} /* (0, 12, 2) {real, imag} */,
  {32'h4405d1ff, 32'h42fee4dc} /* (0, 12, 1) {real, imag} */,
  {32'h4365b1bc, 32'h00000000} /* (0, 12, 0) {real, imag} */,
  {32'h43c56c44, 32'hc2733e44} /* (0, 11, 31) {real, imag} */,
  {32'hc36695ef, 32'h42b2079e} /* (0, 11, 30) {real, imag} */,
  {32'hc16fa73c, 32'hc14459a4} /* (0, 11, 29) {real, imag} */,
  {32'hc1ed9a5e, 32'hc315a451} /* (0, 11, 28) {real, imag} */,
  {32'hc0975228, 32'h412c3710} /* (0, 11, 27) {real, imag} */,
  {32'h40a4f898, 32'hc0e2c6fc} /* (0, 11, 26) {real, imag} */,
  {32'h3e285b40, 32'h42236a8e} /* (0, 11, 25) {real, imag} */,
  {32'h4177313b, 32'h41408494} /* (0, 11, 24) {real, imag} */,
  {32'h41ad0341, 32'h42209e2c} /* (0, 11, 23) {real, imag} */,
  {32'hc2493922, 32'hc2b7d0f0} /* (0, 11, 22) {real, imag} */,
  {32'hc297ba4a, 32'h42b47295} /* (0, 11, 21) {real, imag} */,
  {32'h427f959a, 32'hc23ed354} /* (0, 11, 20) {real, imag} */,
  {32'h418ff65e, 32'hc1c928e6} /* (0, 11, 19) {real, imag} */,
  {32'h41c11e14, 32'h4078b290} /* (0, 11, 18) {real, imag} */,
  {32'hc19bba2d, 32'h41a081a0} /* (0, 11, 17) {real, imag} */,
  {32'hc1b8db17, 32'h00000000} /* (0, 11, 16) {real, imag} */,
  {32'hc19bba2d, 32'hc1a081a0} /* (0, 11, 15) {real, imag} */,
  {32'h41c11e14, 32'hc078b290} /* (0, 11, 14) {real, imag} */,
  {32'h418ff65e, 32'h41c928e6} /* (0, 11, 13) {real, imag} */,
  {32'h427f959a, 32'h423ed354} /* (0, 11, 12) {real, imag} */,
  {32'hc297ba4a, 32'hc2b47295} /* (0, 11, 11) {real, imag} */,
  {32'hc2493922, 32'h42b7d0f0} /* (0, 11, 10) {real, imag} */,
  {32'h41ad0341, 32'hc2209e2c} /* (0, 11, 9) {real, imag} */,
  {32'h4177313b, 32'hc1408494} /* (0, 11, 8) {real, imag} */,
  {32'h3e285b40, 32'hc2236a8e} /* (0, 11, 7) {real, imag} */,
  {32'h40a4f898, 32'h40e2c6fc} /* (0, 11, 6) {real, imag} */,
  {32'hc0975228, 32'hc12c3710} /* (0, 11, 5) {real, imag} */,
  {32'hc1ed9a5e, 32'h4315a451} /* (0, 11, 4) {real, imag} */,
  {32'hc16fa73c, 32'h414459a4} /* (0, 11, 3) {real, imag} */,
  {32'hc36695ef, 32'hc2b2079e} /* (0, 11, 2) {real, imag} */,
  {32'h43c56c44, 32'h42733e44} /* (0, 11, 1) {real, imag} */,
  {32'h42208620, 32'h00000000} /* (0, 11, 0) {real, imag} */,
  {32'h426f3904, 32'h42071956} /* (0, 10, 31) {real, imag} */,
  {32'h42d8c5ea, 32'h42aede09} /* (0, 10, 30) {real, imag} */,
  {32'hc2852448, 32'hc273bd8f} /* (0, 10, 29) {real, imag} */,
  {32'hc212f00a, 32'hc1931898} /* (0, 10, 28) {real, imag} */,
  {32'h426ca2ae, 32'hc299dfce} /* (0, 10, 27) {real, imag} */,
  {32'hc2478ece, 32'hc1e1b279} /* (0, 10, 26) {real, imag} */,
  {32'hc1c77988, 32'h42a4c536} /* (0, 10, 25) {real, imag} */,
  {32'h42d178ac, 32'hc13d756e} /* (0, 10, 24) {real, imag} */,
  {32'h422ba17e, 32'hc1899d3c} /* (0, 10, 23) {real, imag} */,
  {32'h42ea34b8, 32'h413982aa} /* (0, 10, 22) {real, imag} */,
  {32'h41160a4e, 32'hc2784646} /* (0, 10, 21) {real, imag} */,
  {32'hc1966992, 32'h4245ec58} /* (0, 10, 20) {real, imag} */,
  {32'hbfeb0d68, 32'hc1a22146} /* (0, 10, 19) {real, imag} */,
  {32'hc2cda4c7, 32'hc23eff91} /* (0, 10, 18) {real, imag} */,
  {32'hc1978cfa, 32'h403cc840} /* (0, 10, 17) {real, imag} */,
  {32'h42c2355b, 32'h00000000} /* (0, 10, 16) {real, imag} */,
  {32'hc1978cfa, 32'hc03cc840} /* (0, 10, 15) {real, imag} */,
  {32'hc2cda4c7, 32'h423eff91} /* (0, 10, 14) {real, imag} */,
  {32'hbfeb0d68, 32'h41a22146} /* (0, 10, 13) {real, imag} */,
  {32'hc1966992, 32'hc245ec58} /* (0, 10, 12) {real, imag} */,
  {32'h41160a4e, 32'h42784646} /* (0, 10, 11) {real, imag} */,
  {32'h42ea34b8, 32'hc13982aa} /* (0, 10, 10) {real, imag} */,
  {32'h422ba17e, 32'h41899d3c} /* (0, 10, 9) {real, imag} */,
  {32'h42d178ac, 32'h413d756e} /* (0, 10, 8) {real, imag} */,
  {32'hc1c77988, 32'hc2a4c536} /* (0, 10, 7) {real, imag} */,
  {32'hc2478ece, 32'h41e1b279} /* (0, 10, 6) {real, imag} */,
  {32'h426ca2ae, 32'h4299dfce} /* (0, 10, 5) {real, imag} */,
  {32'hc212f00a, 32'h41931898} /* (0, 10, 4) {real, imag} */,
  {32'hc2852448, 32'h4273bd8f} /* (0, 10, 3) {real, imag} */,
  {32'h42d8c5ea, 32'hc2aede09} /* (0, 10, 2) {real, imag} */,
  {32'h426f3904, 32'hc2071956} /* (0, 10, 1) {real, imag} */,
  {32'hc395ee72, 32'h00000000} /* (0, 10, 0) {real, imag} */,
  {32'hc3328cb8, 32'h43173d1a} /* (0, 9, 31) {real, imag} */,
  {32'h4310dd07, 32'hc1ab9f16} /* (0, 9, 30) {real, imag} */,
  {32'h3ec7b500, 32'h401c0a18} /* (0, 9, 29) {real, imag} */,
  {32'hc239e70f, 32'h426d0f3e} /* (0, 9, 28) {real, imag} */,
  {32'h42335af7, 32'hc3002be2} /* (0, 9, 27) {real, imag} */,
  {32'hc1f961b4, 32'h41a87cc6} /* (0, 9, 26) {real, imag} */,
  {32'hc23f8e45, 32'h413173c4} /* (0, 9, 25) {real, imag} */,
  {32'h421e7296, 32'hc224917c} /* (0, 9, 24) {real, imag} */,
  {32'hbe9d6540, 32'hc18f731d} /* (0, 9, 23) {real, imag} */,
  {32'hc20c636a, 32'hc1ade4be} /* (0, 9, 22) {real, imag} */,
  {32'h42bb8a76, 32'hc246a202} /* (0, 9, 21) {real, imag} */,
  {32'h41c8fa21, 32'h41694884} /* (0, 9, 20) {real, imag} */,
  {32'hc27a0bf0, 32'hc11b369f} /* (0, 9, 19) {real, imag} */,
  {32'h423d11ef, 32'hbdd96700} /* (0, 9, 18) {real, imag} */,
  {32'hc1832db0, 32'hc21f4e38} /* (0, 9, 17) {real, imag} */,
  {32'h40545210, 32'h00000000} /* (0, 9, 16) {real, imag} */,
  {32'hc1832db0, 32'h421f4e38} /* (0, 9, 15) {real, imag} */,
  {32'h423d11ef, 32'h3dd96700} /* (0, 9, 14) {real, imag} */,
  {32'hc27a0bf0, 32'h411b369f} /* (0, 9, 13) {real, imag} */,
  {32'h41c8fa21, 32'hc1694884} /* (0, 9, 12) {real, imag} */,
  {32'h42bb8a76, 32'h4246a202} /* (0, 9, 11) {real, imag} */,
  {32'hc20c636a, 32'h41ade4be} /* (0, 9, 10) {real, imag} */,
  {32'hbe9d6540, 32'h418f731d} /* (0, 9, 9) {real, imag} */,
  {32'h421e7296, 32'h4224917c} /* (0, 9, 8) {real, imag} */,
  {32'hc23f8e45, 32'hc13173c4} /* (0, 9, 7) {real, imag} */,
  {32'hc1f961b4, 32'hc1a87cc6} /* (0, 9, 6) {real, imag} */,
  {32'h42335af7, 32'h43002be2} /* (0, 9, 5) {real, imag} */,
  {32'hc239e70f, 32'hc26d0f3e} /* (0, 9, 4) {real, imag} */,
  {32'h3ec7b500, 32'hc01c0a18} /* (0, 9, 3) {real, imag} */,
  {32'h4310dd07, 32'h41ab9f16} /* (0, 9, 2) {real, imag} */,
  {32'hc3328cb8, 32'hc3173d1a} /* (0, 9, 1) {real, imag} */,
  {32'hc3b681ee, 32'h00000000} /* (0, 9, 0) {real, imag} */,
  {32'hc399c9a0, 32'h436368c3} /* (0, 8, 31) {real, imag} */,
  {32'h4358b519, 32'hc0b75240} /* (0, 8, 30) {real, imag} */,
  {32'hc232ffc5, 32'hc285e444} /* (0, 8, 29) {real, imag} */,
  {32'hc23d2488, 32'hc24e1e18} /* (0, 8, 28) {real, imag} */,
  {32'h4244d291, 32'hc1ecff0a} /* (0, 8, 27) {real, imag} */,
  {32'hc18324b4, 32'hc28c3a13} /* (0, 8, 26) {real, imag} */,
  {32'hc1f94048, 32'h40a75aec} /* (0, 8, 25) {real, imag} */,
  {32'h4205b75b, 32'hc25120d3} /* (0, 8, 24) {real, imag} */,
  {32'hc0e78a50, 32'h40e4a640} /* (0, 8, 23) {real, imag} */,
  {32'hc235222a, 32'hc0a06848} /* (0, 8, 22) {real, imag} */,
  {32'h405f2d40, 32'h41c1e599} /* (0, 8, 21) {real, imag} */,
  {32'hc11b6a62, 32'hc14d33e1} /* (0, 8, 20) {real, imag} */,
  {32'h41fd7255, 32'h41a6cd89} /* (0, 8, 19) {real, imag} */,
  {32'h40ea1f2c, 32'h405ad660} /* (0, 8, 18) {real, imag} */,
  {32'hc101751e, 32'hc20ac3f7} /* (0, 8, 17) {real, imag} */,
  {32'hc10dd17b, 32'h00000000} /* (0, 8, 16) {real, imag} */,
  {32'hc101751e, 32'h420ac3f7} /* (0, 8, 15) {real, imag} */,
  {32'h40ea1f2c, 32'hc05ad660} /* (0, 8, 14) {real, imag} */,
  {32'h41fd7255, 32'hc1a6cd89} /* (0, 8, 13) {real, imag} */,
  {32'hc11b6a62, 32'h414d33e1} /* (0, 8, 12) {real, imag} */,
  {32'h405f2d40, 32'hc1c1e599} /* (0, 8, 11) {real, imag} */,
  {32'hc235222a, 32'h40a06848} /* (0, 8, 10) {real, imag} */,
  {32'hc0e78a50, 32'hc0e4a640} /* (0, 8, 9) {real, imag} */,
  {32'h4205b75b, 32'h425120d3} /* (0, 8, 8) {real, imag} */,
  {32'hc1f94048, 32'hc0a75aec} /* (0, 8, 7) {real, imag} */,
  {32'hc18324b4, 32'h428c3a13} /* (0, 8, 6) {real, imag} */,
  {32'h4244d291, 32'h41ecff0a} /* (0, 8, 5) {real, imag} */,
  {32'hc23d2488, 32'h424e1e18} /* (0, 8, 4) {real, imag} */,
  {32'hc232ffc5, 32'h4285e444} /* (0, 8, 3) {real, imag} */,
  {32'h4358b519, 32'h40b75240} /* (0, 8, 2) {real, imag} */,
  {32'hc399c9a0, 32'hc36368c3} /* (0, 8, 1) {real, imag} */,
  {32'hc3b2bb57, 32'h00000000} /* (0, 8, 0) {real, imag} */,
  {32'hc3d95da4, 32'h434252e2} /* (0, 7, 31) {real, imag} */,
  {32'h437a708e, 32'h419bd0e8} /* (0, 7, 30) {real, imag} */,
  {32'h40e01550, 32'hc1c2524c} /* (0, 7, 29) {real, imag} */,
  {32'hc27a416f, 32'hc2e3c718} /* (0, 7, 28) {real, imag} */,
  {32'h42afc4c4, 32'h42735e6b} /* (0, 7, 27) {real, imag} */,
  {32'hc28c6170, 32'hc280ec00} /* (0, 7, 26) {real, imag} */,
  {32'h41cf35dd, 32'hc26da2ec} /* (0, 7, 25) {real, imag} */,
  {32'h4288e301, 32'hc20c8238} /* (0, 7, 24) {real, imag} */,
  {32'h426e8e9a, 32'h42103279} /* (0, 7, 23) {real, imag} */,
  {32'h4135fb43, 32'hc081be00} /* (0, 7, 22) {real, imag} */,
  {32'h42270d86, 32'hc17b2c58} /* (0, 7, 21) {real, imag} */,
  {32'h420cfcf5, 32'h428ed8dc} /* (0, 7, 20) {real, imag} */,
  {32'h421016ca, 32'hc2668ce7} /* (0, 7, 19) {real, imag} */,
  {32'h41a673a3, 32'hc0975c26} /* (0, 7, 18) {real, imag} */,
  {32'h3f84c4e0, 32'h4196621a} /* (0, 7, 17) {real, imag} */,
  {32'h4196b696, 32'h00000000} /* (0, 7, 16) {real, imag} */,
  {32'h3f84c4e0, 32'hc196621a} /* (0, 7, 15) {real, imag} */,
  {32'h41a673a3, 32'h40975c26} /* (0, 7, 14) {real, imag} */,
  {32'h421016ca, 32'h42668ce7} /* (0, 7, 13) {real, imag} */,
  {32'h420cfcf5, 32'hc28ed8dc} /* (0, 7, 12) {real, imag} */,
  {32'h42270d86, 32'h417b2c58} /* (0, 7, 11) {real, imag} */,
  {32'h4135fb43, 32'h4081be00} /* (0, 7, 10) {real, imag} */,
  {32'h426e8e9a, 32'hc2103279} /* (0, 7, 9) {real, imag} */,
  {32'h4288e301, 32'h420c8238} /* (0, 7, 8) {real, imag} */,
  {32'h41cf35dd, 32'h426da2ec} /* (0, 7, 7) {real, imag} */,
  {32'hc28c6170, 32'h4280ec00} /* (0, 7, 6) {real, imag} */,
  {32'h42afc4c4, 32'hc2735e6b} /* (0, 7, 5) {real, imag} */,
  {32'hc27a416f, 32'h42e3c718} /* (0, 7, 4) {real, imag} */,
  {32'h40e01550, 32'h41c2524c} /* (0, 7, 3) {real, imag} */,
  {32'h437a708e, 32'hc19bd0e8} /* (0, 7, 2) {real, imag} */,
  {32'hc3d95da4, 32'hc34252e2} /* (0, 7, 1) {real, imag} */,
  {32'hc3e4a1ff, 32'h00000000} /* (0, 7, 0) {real, imag} */,
  {32'hc3c39e14, 32'h4384d214} /* (0, 6, 31) {real, imag} */,
  {32'h43b0ed1e, 32'h42c8de3b} /* (0, 6, 30) {real, imag} */,
  {32'h42b20232, 32'hc1f46dee} /* (0, 6, 29) {real, imag} */,
  {32'hc2b12354, 32'hc1a9b674} /* (0, 6, 28) {real, imag} */,
  {32'h42ad97ea, 32'h411f27f4} /* (0, 6, 27) {real, imag} */,
  {32'hc1d417f9, 32'hc2115142} /* (0, 6, 26) {real, imag} */,
  {32'hc208a6f6, 32'h42193832} /* (0, 6, 25) {real, imag} */,
  {32'hc03356a0, 32'hc2756198} /* (0, 6, 24) {real, imag} */,
  {32'h418ecd7c, 32'hc11e9a26} /* (0, 6, 23) {real, imag} */,
  {32'hc1bce11e, 32'h42f9a577} /* (0, 6, 22) {real, imag} */,
  {32'h428d86d0, 32'hc1dbaca2} /* (0, 6, 21) {real, imag} */,
  {32'hc284123a, 32'h41cec01c} /* (0, 6, 20) {real, imag} */,
  {32'h42301b92, 32'h421dc658} /* (0, 6, 19) {real, imag} */,
  {32'h4266d4a0, 32'h406f965e} /* (0, 6, 18) {real, imag} */,
  {32'hc2207ada, 32'hc215445a} /* (0, 6, 17) {real, imag} */,
  {32'hc2233935, 32'h00000000} /* (0, 6, 16) {real, imag} */,
  {32'hc2207ada, 32'h4215445a} /* (0, 6, 15) {real, imag} */,
  {32'h4266d4a0, 32'hc06f965e} /* (0, 6, 14) {real, imag} */,
  {32'h42301b92, 32'hc21dc658} /* (0, 6, 13) {real, imag} */,
  {32'hc284123a, 32'hc1cec01c} /* (0, 6, 12) {real, imag} */,
  {32'h428d86d0, 32'h41dbaca2} /* (0, 6, 11) {real, imag} */,
  {32'hc1bce11e, 32'hc2f9a577} /* (0, 6, 10) {real, imag} */,
  {32'h418ecd7c, 32'h411e9a26} /* (0, 6, 9) {real, imag} */,
  {32'hc03356a0, 32'h42756198} /* (0, 6, 8) {real, imag} */,
  {32'hc208a6f6, 32'hc2193832} /* (0, 6, 7) {real, imag} */,
  {32'hc1d417f9, 32'h42115142} /* (0, 6, 6) {real, imag} */,
  {32'h42ad97ea, 32'hc11f27f4} /* (0, 6, 5) {real, imag} */,
  {32'hc2b12354, 32'h41a9b674} /* (0, 6, 4) {real, imag} */,
  {32'h42b20232, 32'h41f46dee} /* (0, 6, 3) {real, imag} */,
  {32'h43b0ed1e, 32'hc2c8de3b} /* (0, 6, 2) {real, imag} */,
  {32'hc3c39e14, 32'hc384d214} /* (0, 6, 1) {real, imag} */,
  {32'hc407327b, 32'h00000000} /* (0, 6, 0) {real, imag} */,
  {32'hc38feea2, 32'h43f730f0} /* (0, 5, 31) {real, imag} */,
  {32'h42361de8, 32'h42b4c4c0} /* (0, 5, 30) {real, imag} */,
  {32'h42eec432, 32'h40be72f8} /* (0, 5, 29) {real, imag} */,
  {32'hc19417f6, 32'hc19c4000} /* (0, 5, 28) {real, imag} */,
  {32'h42cdaccd, 32'h41920572} /* (0, 5, 27) {real, imag} */,
  {32'hc22a187f, 32'hc2ceb9bc} /* (0, 5, 26) {real, imag} */,
  {32'h412df3b8, 32'hc1f9d8ca} /* (0, 5, 25) {real, imag} */,
  {32'hc1e686e6, 32'h41d55cab} /* (0, 5, 24) {real, imag} */,
  {32'h425b052b, 32'h42ad5d4a} /* (0, 5, 23) {real, imag} */,
  {32'h41b8c385, 32'hc14d5ff8} /* (0, 5, 22) {real, imag} */,
  {32'h4032eb78, 32'hc21d60d3} /* (0, 5, 21) {real, imag} */,
  {32'h428e9720, 32'hc2705738} /* (0, 5, 20) {real, imag} */,
  {32'h40e1ae56, 32'hc1b8a10e} /* (0, 5, 19) {real, imag} */,
  {32'h42076219, 32'h41e10fd6} /* (0, 5, 18) {real, imag} */,
  {32'hc110cc82, 32'h402cb040} /* (0, 5, 17) {real, imag} */,
  {32'h42801440, 32'h00000000} /* (0, 5, 16) {real, imag} */,
  {32'hc110cc82, 32'hc02cb040} /* (0, 5, 15) {real, imag} */,
  {32'h42076219, 32'hc1e10fd6} /* (0, 5, 14) {real, imag} */,
  {32'h40e1ae56, 32'h41b8a10e} /* (0, 5, 13) {real, imag} */,
  {32'h428e9720, 32'h42705738} /* (0, 5, 12) {real, imag} */,
  {32'h4032eb78, 32'h421d60d3} /* (0, 5, 11) {real, imag} */,
  {32'h41b8c385, 32'h414d5ff8} /* (0, 5, 10) {real, imag} */,
  {32'h425b052b, 32'hc2ad5d4a} /* (0, 5, 9) {real, imag} */,
  {32'hc1e686e6, 32'hc1d55cab} /* (0, 5, 8) {real, imag} */,
  {32'h412df3b8, 32'h41f9d8ca} /* (0, 5, 7) {real, imag} */,
  {32'hc22a187f, 32'h42ceb9bc} /* (0, 5, 6) {real, imag} */,
  {32'h42cdaccd, 32'hc1920572} /* (0, 5, 5) {real, imag} */,
  {32'hc19417f6, 32'h419c4000} /* (0, 5, 4) {real, imag} */,
  {32'h42eec432, 32'hc0be72f8} /* (0, 5, 3) {real, imag} */,
  {32'h42361de8, 32'hc2b4c4c0} /* (0, 5, 2) {real, imag} */,
  {32'hc38feea2, 32'hc3f730f0} /* (0, 5, 1) {real, imag} */,
  {32'hc45143bc, 32'h00000000} /* (0, 5, 0) {real, imag} */,
  {32'hc3973c29, 32'h441b355f} /* (0, 4, 31) {real, imag} */,
  {32'hc2e6090a, 32'hc1ffde1e} /* (0, 4, 30) {real, imag} */,
  {32'h42ba47e8, 32'h42461bcf} /* (0, 4, 29) {real, imag} */,
  {32'h42582505, 32'hc2e57123} /* (0, 4, 28) {real, imag} */,
  {32'h42aa81e6, 32'h42a55a43} /* (0, 4, 27) {real, imag} */,
  {32'hc18cb7a0, 32'hc2ac4c22} /* (0, 4, 26) {real, imag} */,
  {32'hbc4c2c00, 32'hc1356755} /* (0, 4, 25) {real, imag} */,
  {32'hc2ccbed6, 32'h3fc7a340} /* (0, 4, 24) {real, imag} */,
  {32'h42c175aa, 32'hc10722d6} /* (0, 4, 23) {real, imag} */,
  {32'hc1fcc1f5, 32'h41859eda} /* (0, 4, 22) {real, imag} */,
  {32'h42e34640, 32'h4231d8b4} /* (0, 4, 21) {real, imag} */,
  {32'hc1a05e9e, 32'h41667dd8} /* (0, 4, 20) {real, imag} */,
  {32'h40ff31f8, 32'hbee93e00} /* (0, 4, 19) {real, imag} */,
  {32'h427ea882, 32'hc29dd3db} /* (0, 4, 18) {real, imag} */,
  {32'hc09d164d, 32'hc1f4ac3b} /* (0, 4, 17) {real, imag} */,
  {32'hc1e0631a, 32'h00000000} /* (0, 4, 16) {real, imag} */,
  {32'hc09d164d, 32'h41f4ac3b} /* (0, 4, 15) {real, imag} */,
  {32'h427ea882, 32'h429dd3db} /* (0, 4, 14) {real, imag} */,
  {32'h40ff31f8, 32'h3ee93e00} /* (0, 4, 13) {real, imag} */,
  {32'hc1a05e9e, 32'hc1667dd8} /* (0, 4, 12) {real, imag} */,
  {32'h42e34640, 32'hc231d8b4} /* (0, 4, 11) {real, imag} */,
  {32'hc1fcc1f5, 32'hc1859eda} /* (0, 4, 10) {real, imag} */,
  {32'h42c175aa, 32'h410722d6} /* (0, 4, 9) {real, imag} */,
  {32'hc2ccbed6, 32'hbfc7a340} /* (0, 4, 8) {real, imag} */,
  {32'hbc4c2c00, 32'h41356755} /* (0, 4, 7) {real, imag} */,
  {32'hc18cb7a0, 32'h42ac4c22} /* (0, 4, 6) {real, imag} */,
  {32'h42aa81e6, 32'hc2a55a43} /* (0, 4, 5) {real, imag} */,
  {32'h42582505, 32'h42e57123} /* (0, 4, 4) {real, imag} */,
  {32'h42ba47e8, 32'hc2461bcf} /* (0, 4, 3) {real, imag} */,
  {32'hc2e6090a, 32'h41ffde1e} /* (0, 4, 2) {real, imag} */,
  {32'hc3973c29, 32'hc41b355f} /* (0, 4, 1) {real, imag} */,
  {32'hc438b5b0, 32'h00000000} /* (0, 4, 0) {real, imag} */,
  {32'hc374df4b, 32'h441edb82} /* (0, 3, 31) {real, imag} */,
  {32'hc2a0216d, 32'hc3414ad2} /* (0, 3, 30) {real, imag} */,
  {32'h42e36777, 32'h41c20278} /* (0, 3, 29) {real, imag} */,
  {32'hc2bd3ea3, 32'hc31d38a0} /* (0, 3, 28) {real, imag} */,
  {32'h429a4f81, 32'h42c5eb6e} /* (0, 3, 27) {real, imag} */,
  {32'h4255ef14, 32'hc194666f} /* (0, 3, 26) {real, imag} */,
  {32'hc1b526aa, 32'hc0db72a0} /* (0, 3, 25) {real, imag} */,
  {32'h3fd15620, 32'hc1a08f65} /* (0, 3, 24) {real, imag} */,
  {32'hc0c535ae, 32'h419c0590} /* (0, 3, 23) {real, imag} */,
  {32'h41789ea6, 32'h41ed1f54} /* (0, 3, 22) {real, imag} */,
  {32'h423b9708, 32'hc21d4bf4} /* (0, 3, 21) {real, imag} */,
  {32'h419a6544, 32'hc174f320} /* (0, 3, 20) {real, imag} */,
  {32'h41f523f2, 32'hc2041ce0} /* (0, 3, 19) {real, imag} */,
  {32'h418579e2, 32'h4202e222} /* (0, 3, 18) {real, imag} */,
  {32'h40315c6c, 32'hc1ff2680} /* (0, 3, 17) {real, imag} */,
  {32'hc1a162f3, 32'h00000000} /* (0, 3, 16) {real, imag} */,
  {32'h40315c6c, 32'h41ff2680} /* (0, 3, 15) {real, imag} */,
  {32'h418579e2, 32'hc202e222} /* (0, 3, 14) {real, imag} */,
  {32'h41f523f2, 32'h42041ce0} /* (0, 3, 13) {real, imag} */,
  {32'h419a6544, 32'h4174f320} /* (0, 3, 12) {real, imag} */,
  {32'h423b9708, 32'h421d4bf4} /* (0, 3, 11) {real, imag} */,
  {32'h41789ea6, 32'hc1ed1f54} /* (0, 3, 10) {real, imag} */,
  {32'hc0c535ae, 32'hc19c0590} /* (0, 3, 9) {real, imag} */,
  {32'h3fd15620, 32'h41a08f65} /* (0, 3, 8) {real, imag} */,
  {32'hc1b526aa, 32'h40db72a0} /* (0, 3, 7) {real, imag} */,
  {32'h4255ef14, 32'h4194666f} /* (0, 3, 6) {real, imag} */,
  {32'h429a4f81, 32'hc2c5eb6e} /* (0, 3, 5) {real, imag} */,
  {32'hc2bd3ea3, 32'h431d38a0} /* (0, 3, 4) {real, imag} */,
  {32'h42e36777, 32'hc1c20278} /* (0, 3, 3) {real, imag} */,
  {32'hc2a0216d, 32'h43414ad2} /* (0, 3, 2) {real, imag} */,
  {32'hc374df4b, 32'hc41edb82} /* (0, 3, 1) {real, imag} */,
  {32'hc435cbf0, 32'h00000000} /* (0, 3, 0) {real, imag} */,
  {32'hc393601c, 32'h440893be} /* (0, 2, 31) {real, imag} */,
  {32'hc338e96b, 32'hc33a2778} /* (0, 2, 30) {real, imag} */,
  {32'h433799cc, 32'h420f5f63} /* (0, 2, 29) {real, imag} */,
  {32'hc2aaceac, 32'hc2b51238} /* (0, 2, 28) {real, imag} */,
  {32'h424bd838, 32'h42956507} /* (0, 2, 27) {real, imag} */,
  {32'hbed34f80, 32'h41194974} /* (0, 2, 26) {real, imag} */,
  {32'hc269b9f0, 32'h42c7db0f} /* (0, 2, 25) {real, imag} */,
  {32'hc0417a98, 32'h4182bc84} /* (0, 2, 24) {real, imag} */,
  {32'h41f007b4, 32'hc228ecf1} /* (0, 2, 23) {real, imag} */,
  {32'hc19e0558, 32'h416e0990} /* (0, 2, 22) {real, imag} */,
  {32'hc0745ff0, 32'hc167cd70} /* (0, 2, 21) {real, imag} */,
  {32'h41bdcc2e, 32'h41858286} /* (0, 2, 20) {real, imag} */,
  {32'hc2318da0, 32'h422332b6} /* (0, 2, 19) {real, imag} */,
  {32'hc1cc2006, 32'h41d41492} /* (0, 2, 18) {real, imag} */,
  {32'h4200aa96, 32'h4110172c} /* (0, 2, 17) {real, imag} */,
  {32'hc1db4f51, 32'h00000000} /* (0, 2, 16) {real, imag} */,
  {32'h4200aa96, 32'hc110172c} /* (0, 2, 15) {real, imag} */,
  {32'hc1cc2006, 32'hc1d41492} /* (0, 2, 14) {real, imag} */,
  {32'hc2318da0, 32'hc22332b6} /* (0, 2, 13) {real, imag} */,
  {32'h41bdcc2e, 32'hc1858286} /* (0, 2, 12) {real, imag} */,
  {32'hc0745ff0, 32'h4167cd70} /* (0, 2, 11) {real, imag} */,
  {32'hc19e0558, 32'hc16e0990} /* (0, 2, 10) {real, imag} */,
  {32'h41f007b4, 32'h4228ecf1} /* (0, 2, 9) {real, imag} */,
  {32'hc0417a98, 32'hc182bc84} /* (0, 2, 8) {real, imag} */,
  {32'hc269b9f0, 32'hc2c7db0f} /* (0, 2, 7) {real, imag} */,
  {32'hbed34f80, 32'hc1194974} /* (0, 2, 6) {real, imag} */,
  {32'h424bd838, 32'hc2956507} /* (0, 2, 5) {real, imag} */,
  {32'hc2aaceac, 32'h42b51238} /* (0, 2, 4) {real, imag} */,
  {32'h433799cc, 32'hc20f5f63} /* (0, 2, 3) {real, imag} */,
  {32'hc338e96b, 32'h433a2778} /* (0, 2, 2) {real, imag} */,
  {32'hc393601c, 32'hc40893be} /* (0, 2, 1) {real, imag} */,
  {32'hc3e75dbd, 32'h00000000} /* (0, 2, 0) {real, imag} */,
  {32'hc3aaab64, 32'h44051d4e} /* (0, 1, 31) {real, imag} */,
  {32'hc394214d, 32'hc330e42e} /* (0, 1, 30) {real, imag} */,
  {32'h431871ed, 32'hc26d5f25} /* (0, 1, 29) {real, imag} */,
  {32'h42401d3b, 32'hc2e1d84b} /* (0, 1, 28) {real, imag} */,
  {32'h4307a697, 32'h42933747} /* (0, 1, 27) {real, imag} */,
  {32'hc1a6dc20, 32'h41fb7c9f} /* (0, 1, 26) {real, imag} */,
  {32'hc23f75e7, 32'h42919701} /* (0, 1, 25) {real, imag} */,
  {32'h3fde3b40, 32'hc28cbce1} /* (0, 1, 24) {real, imag} */,
  {32'h42072930, 32'hc0bed78c} /* (0, 1, 23) {real, imag} */,
  {32'hc1f8d176, 32'h42072126} /* (0, 1, 22) {real, imag} */,
  {32'h42602b36, 32'hc07cb512} /* (0, 1, 21) {real, imag} */,
  {32'hc20a73ed, 32'h42441240} /* (0, 1, 20) {real, imag} */,
  {32'hc2828243, 32'hc19e310d} /* (0, 1, 19) {real, imag} */,
  {32'hc22f7255, 32'hc24845a4} /* (0, 1, 18) {real, imag} */,
  {32'h422e61f0, 32'hc236fc0d} /* (0, 1, 17) {real, imag} */,
  {32'h422dd2ab, 32'h00000000} /* (0, 1, 16) {real, imag} */,
  {32'h422e61f0, 32'h4236fc0d} /* (0, 1, 15) {real, imag} */,
  {32'hc22f7255, 32'h424845a4} /* (0, 1, 14) {real, imag} */,
  {32'hc2828243, 32'h419e310d} /* (0, 1, 13) {real, imag} */,
  {32'hc20a73ed, 32'hc2441240} /* (0, 1, 12) {real, imag} */,
  {32'h42602b36, 32'h407cb512} /* (0, 1, 11) {real, imag} */,
  {32'hc1f8d176, 32'hc2072126} /* (0, 1, 10) {real, imag} */,
  {32'h42072930, 32'h40bed78c} /* (0, 1, 9) {real, imag} */,
  {32'h3fde3b40, 32'h428cbce1} /* (0, 1, 8) {real, imag} */,
  {32'hc23f75e7, 32'hc2919701} /* (0, 1, 7) {real, imag} */,
  {32'hc1a6dc20, 32'hc1fb7c9f} /* (0, 1, 6) {real, imag} */,
  {32'h4307a697, 32'hc2933747} /* (0, 1, 5) {real, imag} */,
  {32'h42401d3b, 32'h42e1d84b} /* (0, 1, 4) {real, imag} */,
  {32'h431871ed, 32'h426d5f25} /* (0, 1, 3) {real, imag} */,
  {32'hc394214d, 32'h4330e42e} /* (0, 1, 2) {real, imag} */,
  {32'hc3aaab64, 32'hc4051d4e} /* (0, 1, 1) {real, imag} */,
  {32'hc389dbcb, 32'h00000000} /* (0, 1, 0) {real, imag} */,
  {32'hc3b70e86, 32'h43ab0c49} /* (0, 0, 31) {real, imag} */,
  {32'hc30917e2, 32'hc2580336} /* (0, 0, 30) {real, imag} */,
  {32'h4277f3d7, 32'h42210366} /* (0, 0, 29) {real, imag} */,
  {32'h423ca4e4, 32'hc29538dd} /* (0, 0, 28) {real, imag} */,
  {32'h4301daf9, 32'h41f04d7e} /* (0, 0, 27) {real, imag} */,
  {32'hc182e4a6, 32'h41251c9b} /* (0, 0, 26) {real, imag} */,
  {32'h420e55d6, 32'h41b1a050} /* (0, 0, 25) {real, imag} */,
  {32'h412a9dba, 32'hc0782400} /* (0, 0, 24) {real, imag} */,
  {32'h42517b5a, 32'hc03c65d0} /* (0, 0, 23) {real, imag} */,
  {32'hc25d6380, 32'hc1b9e944} /* (0, 0, 22) {real, imag} */,
  {32'h41180d26, 32'hc1e228d1} /* (0, 0, 21) {real, imag} */,
  {32'hc1ba4f48, 32'h41ba516d} /* (0, 0, 20) {real, imag} */,
  {32'h4209db67, 32'h426b51e4} /* (0, 0, 19) {real, imag} */,
  {32'hc196b7a5, 32'h422bda54} /* (0, 0, 18) {real, imag} */,
  {32'h410f4220, 32'h4026c440} /* (0, 0, 17) {real, imag} */,
  {32'h41479af4, 32'h00000000} /* (0, 0, 16) {real, imag} */,
  {32'h410f4220, 32'hc026c440} /* (0, 0, 15) {real, imag} */,
  {32'hc196b7a5, 32'hc22bda54} /* (0, 0, 14) {real, imag} */,
  {32'h4209db67, 32'hc26b51e4} /* (0, 0, 13) {real, imag} */,
  {32'hc1ba4f48, 32'hc1ba516d} /* (0, 0, 12) {real, imag} */,
  {32'h41180d26, 32'h41e228d1} /* (0, 0, 11) {real, imag} */,
  {32'hc25d6380, 32'h41b9e944} /* (0, 0, 10) {real, imag} */,
  {32'h42517b5a, 32'h403c65d0} /* (0, 0, 9) {real, imag} */,
  {32'h412a9dba, 32'h40782400} /* (0, 0, 8) {real, imag} */,
  {32'h420e55d6, 32'hc1b1a050} /* (0, 0, 7) {real, imag} */,
  {32'hc182e4a6, 32'hc1251c9b} /* (0, 0, 6) {real, imag} */,
  {32'h4301daf9, 32'hc1f04d7e} /* (0, 0, 5) {real, imag} */,
  {32'h423ca4e4, 32'h429538dd} /* (0, 0, 4) {real, imag} */,
  {32'h4277f3d7, 32'hc2210366} /* (0, 0, 3) {real, imag} */,
  {32'hc30917e2, 32'h42580336} /* (0, 0, 2) {real, imag} */,
  {32'hc3b70e86, 32'hc3ab0c49} /* (0, 0, 1) {real, imag} */,
  {32'hc372fd9b, 32'h00000000} /* (0, 0, 0) {real, imag} */};
